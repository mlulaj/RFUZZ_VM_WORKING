`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module DUT(
  input         clock,
  input         reset,
  input         io_meta_reset,
  input  [34:0] io_inputs,
  output        io_coverage_0,
  output        io_coverage_1,
  output        io_coverage_2,
  output        io_coverage_3,
  output        io_coverage_4,
  output        io_coverage_5,
  output        io_coverage_6,
  output        io_coverage_7,
  output        io_coverage_8,
  output        io_coverage_9,
  output        io_coverage_10,
  output        io_coverage_11,
  output        io_coverage_12,
  output        io_coverage_13,
  output        io_coverage_14,
  output        io_coverage_15,
  output        io_coverage_16,
  output        io_coverage_17,
  output        io_coverage_18,
  output        io_coverage_19,
  output        io_coverage_20,
  output        io_coverage_21,
  output        io_coverage_22,
  output        io_coverage_23,
  output        io_coverage_24,
  output        io_coverage_25,
  output        io_coverage_26,
  output        io_coverage_27,
  output        io_coverage_28,
  output        io_coverage_29,
  output        io_coverage_30,
  output        io_coverage_31,
  output        io_coverage_32,
  output        io_coverage_33,
  output        io_coverage_34,
  output        io_coverage_35,
  output        io_coverage_36,
  output        io_coverage_37,
  output        io_coverage_38,
  output        io_coverage_39,
  output        io_coverage_40,
  output        io_coverage_41,
  output        io_coverage_42,
  output        io_coverage_43,
  output        io_coverage_44,
  output        io_coverage_45,
  output        io_coverage_46,
  output        io_coverage_47,
  output        io_coverage_48,
  output        io_coverage_49,
  output        io_coverage_50,
  output        io_coverage_51,
  output        io_coverage_52,
  output        io_coverage_53,
  output        io_coverage_54,
  output        io_coverage_55,
  output        io_coverage_56,
  output        io_coverage_57,
  output        io_coverage_58,
  output        io_coverage_59,
  output        io_coverage_60,
  output        io_coverage_61,
  output        io_coverage_62,
  output        io_coverage_63,
  output        io_coverage_64,
  output        io_coverage_65,
  output        io_coverage_66,
  output        io_coverage_67,
  output        io_coverage_68,
  output        io_coverage_69,
  output        io_coverage_70,
  output        io_coverage_71,
  output        io_coverage_72,
  output        io_coverage_73,
  output        io_coverage_74,
  output        io_coverage_75,
  output        io_coverage_76,
  output        io_coverage_77,
  output        io_coverage_78,
  output        io_coverage_79,
  output        io_coverage_80,
  output        io_coverage_81,
  output        io_coverage_82,
  output        io_coverage_83,
  output        io_coverage_84,
  output        io_coverage_85,
  output        io_coverage_86,
  output        io_coverage_87,
  output        io_coverage_88,
  output        io_coverage_89,
  output        io_coverage_90,
  output        io_coverage_91,
  output        io_coverage_92,
  output        io_coverage_93,
  output        io_coverage_94,
  output        io_coverage_95,
  output        io_coverage_96,
  output        io_coverage_97,
  output        io_coverage_98,
  output        io_coverage_99,
  output        io_coverage_100,
  output        io_coverage_101,
  output        io_coverage_102,
  output        io_coverage_103,
  output        io_coverage_104,
  output        io_coverage_105,
  output        io_coverage_106,
  output        io_coverage_107,
  output        io_coverage_108,
  output        io_coverage_109,
  output        io_coverage_110,
  output        io_coverage_111,
  output        io_coverage_112,
  output        io_coverage_113,
  output        io_coverage_114,
  output        io_coverage_115,
  output        io_coverage_116,
  output        io_coverage_117,
  output        io_coverage_118,
  output        io_coverage_119,
  output        io_coverage_120,
  output        io_coverage_121,
  output        io_coverage_122,
  output        io_coverage_123,
  output        io_coverage_124,
  output        io_coverage_125,
  output        io_coverage_126,
  output        io_coverage_127,
  output        io_coverage_128,
  output        io_coverage_129,
  output        io_coverage_130,
  output        io_coverage_131,
  output        io_coverage_132,
  output        io_coverage_133,
  output        io_coverage_134,
  output        io_coverage_135,
  output        io_coverage_136,
  output        io_coverage_137,
  output        io_coverage_138,
  output        io_coverage_139,
  output        io_coverage_140,
  output        io_coverage_141,
  output        io_coverage_142,
  output        io_coverage_143,
  output        io_coverage_144,
  output        io_coverage_145,
  output        io_coverage_146,
  output        io_coverage_147,
  output        io_coverage_148,
  output        io_coverage_149,
  output        io_coverage_150,
  output        io_coverage_151,
  output        io_coverage_152,
  output        io_coverage_153,
  output        io_coverage_154,
  output        io_coverage_155,
  output        io_coverage_156,
  output        io_coverage_157,
  output        io_coverage_158,
  output        io_coverage_159,
  output        io_coverage_160,
  output        io_coverage_161,
  output        io_coverage_162,
  output        io_coverage_163,
  output        io_coverage_164,
  output        io_coverage_165,
  output        io_coverage_166,
  output        io_coverage_167,
  output        io_coverage_168,
  output        io_coverage_169,
  output        io_coverage_170,
  output        io_coverage_171,
  output        io_coverage_172,
  output        io_coverage_173,
  output        io_coverage_174,
  output        io_coverage_175,
  output        io_coverage_176,
  output        io_coverage_177,
  output        io_coverage_178,
  output        io_coverage_179,
  output        io_coverage_180,
  output        io_coverage_181,
  output        io_coverage_182,
  output        io_coverage_183,
  output        io_coverage_184,
  output        io_coverage_185,
  output        io_coverage_186,
  output        io_coverage_187,
  output        io_coverage_188,
  output        io_coverage_189,
  output        io_coverage_190,
  output        io_coverage_191
);
  wire  bb_clock;
  wire  bb_reset;
  wire  bb_metaReset;
  wire [31:0] bb_io_imem_resp_bits_data;
  wire  bb_io_imem_req_ready;
  wire  bb_io_imem_resp_valid;
  wire  bb_io_reset;
  wire  bb_assert_out;
  wire [745:0] bb_auto_cover_out;
  wire [31:0] _T_202;
  wire  _T_203;
  wire  _T_204;
  wire  _T_205;
  wire  coverage_0;
  wire  coverage_1;
  wire  coverage_2;
  wire  coverage_3;
  wire  coverage_4;
  wire  coverage_5;
  wire  coverage_6;
  wire  coverage_7;
  wire  coverage_8;
  wire  coverage_9;
  wire  coverage_10;
  wire  coverage_11;
  wire  coverage_12;
  wire  coverage_13;
  wire  coverage_14;
  wire  coverage_15;
  wire  coverage_16;
  wire  coverage_17;
  wire  coverage_18;
  wire  coverage_19;
  wire  coverage_20;
  wire  coverage_21;
  wire  coverage_22;
  wire  coverage_23;
  wire  coverage_24;
  wire  coverage_25;
  wire  coverage_26;
  wire  coverage_27;
  wire  coverage_28;
  wire  coverage_29;
  wire  coverage_30;
  wire  coverage_31;
  wire  coverage_32;
  wire  coverage_33;
  wire  coverage_34;
  wire  coverage_35;
  wire  coverage_36;
  wire  coverage_37;
  wire  coverage_38;
  wire  coverage_39;
  wire  coverage_40;
  wire  coverage_41;
  wire  coverage_42;
  wire  coverage_43;
  wire  coverage_44;
  wire  coverage_45;
  wire  coverage_46;
  wire  coverage_47;
  wire  coverage_48;
  wire  coverage_49;
  wire  coverage_50;
  wire  coverage_51;
  wire  coverage_52;
  wire  coverage_53;
  wire  coverage_54;
  wire  coverage_55;
  wire  coverage_56;
  wire  coverage_57;
  wire  coverage_58;
  wire  coverage_59;
  wire  coverage_60;
  wire  coverage_61;
  wire  coverage_62;
  wire  coverage_63;
  wire  coverage_64;
  wire  coverage_65;
  wire  coverage_66;
  wire  coverage_67;
  wire  coverage_68;
  wire  coverage_69;
  wire  coverage_70;
  wire  coverage_71;
  wire  coverage_72;
  wire  coverage_73;
  wire  coverage_74;
  wire  coverage_75;
  wire  coverage_76;
  wire  coverage_77;
  wire  coverage_78;
  wire  coverage_79;
  wire  coverage_80;
  wire  coverage_81;
  wire  coverage_82;
  wire  coverage_83;
  wire  coverage_84;
  wire  coverage_85;
  wire  coverage_86;
  wire  coverage_87;
  wire  coverage_88;
  wire  coverage_89;
  wire  coverage_90;
  wire  coverage_91;
  wire  coverage_92;
  wire  coverage_93;
  wire  coverage_94;
  wire  coverage_95;
  wire  coverage_96;
  wire  coverage_97;
  wire  coverage_98;
  wire  coverage_99;
  wire  coverage_100;
  wire  coverage_101;
  wire  coverage_102;
  wire  coverage_103;
  wire  coverage_104;
  wire  coverage_105;
  wire  coverage_106;
  wire  coverage_107;
  wire  coverage_108;
  wire  coverage_109;
  wire  coverage_110;
  wire  coverage_111;
  wire  coverage_112;
  wire  coverage_113;
  wire  coverage_114;
  wire  coverage_115;
  wire  coverage_116;
  wire  coverage_117;
  wire  coverage_118;
  wire  coverage_119;
  wire  coverage_120;
  wire  coverage_121;
  wire  coverage_122;
  wire  coverage_123;
  wire  coverage_124;
  wire  coverage_125;
  wire  coverage_126;
  wire  coverage_127;
  wire  coverage_128;
  wire  coverage_129;
  wire  coverage_130;
  wire  coverage_131;
  wire  coverage_132;
  wire  coverage_133;
  wire  coverage_134;
  wire  coverage_135;
  wire  coverage_136;
  wire  coverage_137;
  wire  coverage_138;
  wire  coverage_139;
  wire  coverage_140;
  wire  coverage_141;
  wire  coverage_142;
  wire  coverage_143;
  wire  coverage_144;
  wire  coverage_145;
  wire  coverage_146;
  wire  coverage_147;
  wire  coverage_148;
  wire  coverage_149;
  wire  coverage_150;
  wire  coverage_151;
  wire  coverage_152;
  wire  coverage_153;
  wire  coverage_154;
  wire  coverage_155;
  wire  coverage_156;
  wire  coverage_157;
  wire  coverage_158;
  wire  coverage_159;
  wire  coverage_160;
  wire  coverage_161;
  wire  coverage_162;
  wire  coverage_163;
  wire  coverage_164;
  wire  coverage_165;
  wire  coverage_166;
  wire  coverage_167;
  wire  coverage_168;
  wire  coverage_169;
  wire  coverage_170;
  wire  coverage_171;
  wire  coverage_172;
  wire  coverage_173;
  wire  coverage_174;
  wire  coverage_175;
  wire  coverage_176;
  wire  coverage_177;
  wire  coverage_178;
  wire  coverage_179;
  wire  coverage_180;
  wire  coverage_181;
  wire  coverage_182;
  wire  coverage_183;
  wire  coverage_184;
  wire  coverage_185;
  wire  coverage_186;
  wire  coverage_187;
  wire  coverage_188;
  wire  coverage_189;
  wire  coverage_190;
  wire  coverage_191;
  Sodor3Stage bb (
    .clock(bb_clock),
    .reset(bb_reset),
    .metaReset(bb_metaReset),
    .io_imem_resp_bits_data(bb_io_imem_resp_bits_data),
    .io_imem_req_ready(bb_io_imem_req_ready),
    .io_imem_resp_valid(bb_io_imem_resp_valid),
    .io_reset(bb_io_reset),
    .assert_out(bb_assert_out),
    .auto_cover_out(bb_auto_cover_out)
  );
  assign _T_202 = io_inputs[34:3];
  assign _T_203 = io_inputs[2];
  assign _T_204 = io_inputs[1];
  assign _T_205 = io_inputs[0];
  assign coverage_0 = bb_assert_out;
  assign coverage_1 = bb_auto_cover_out[745];
  assign coverage_2 = bb_auto_cover_out[744];
  assign coverage_3 = bb_auto_cover_out[734];
  assign coverage_4 = bb_auto_cover_out[733];
  assign coverage_5 = bb_auto_cover_out[732];
  assign coverage_6 = bb_auto_cover_out[731];
  assign coverage_7 = bb_auto_cover_out[730];
  assign coverage_8 = bb_auto_cover_out[729];
  assign coverage_9 = bb_auto_cover_out[728];
  assign coverage_10 = bb_auto_cover_out[727];
  assign coverage_11 = bb_auto_cover_out[726];
  assign coverage_12 = bb_auto_cover_out[725];
  assign coverage_13 = bb_auto_cover_out[724];
  assign coverage_14 = bb_auto_cover_out[723];
  assign coverage_15 = bb_auto_cover_out[722];
  assign coverage_16 = bb_auto_cover_out[721];
  assign coverage_17 = bb_auto_cover_out[720];
  assign coverage_18 = bb_auto_cover_out[719];
  assign coverage_19 = bb_auto_cover_out[718];
  assign coverage_20 = bb_auto_cover_out[717];
  assign coverage_21 = bb_auto_cover_out[716];
  assign coverage_22 = bb_auto_cover_out[715];
  assign coverage_23 = bb_auto_cover_out[714];
  assign coverage_24 = bb_auto_cover_out[713];
  assign coverage_25 = bb_auto_cover_out[712];
  assign coverage_26 = bb_auto_cover_out[711];
  assign coverage_27 = bb_auto_cover_out[710];
  assign coverage_28 = bb_auto_cover_out[709];
  assign coverage_29 = bb_auto_cover_out[708];
  assign coverage_30 = bb_auto_cover_out[707];
  assign coverage_31 = bb_auto_cover_out[706];
  assign coverage_32 = bb_auto_cover_out[705];
  assign coverage_33 = bb_auto_cover_out[704];
  assign coverage_34 = bb_auto_cover_out[703];
  assign coverage_35 = bb_auto_cover_out[702];
  assign coverage_36 = bb_auto_cover_out[701];
  assign coverage_37 = bb_auto_cover_out[700];
  assign coverage_38 = bb_auto_cover_out[699];
  assign coverage_39 = bb_auto_cover_out[698];
  assign coverage_40 = bb_auto_cover_out[697];
  assign coverage_41 = bb_auto_cover_out[696];
  assign coverage_42 = bb_auto_cover_out[695];
  assign coverage_43 = bb_auto_cover_out[694];
  assign coverage_44 = bb_auto_cover_out[693];
  assign coverage_45 = bb_auto_cover_out[692];
  assign coverage_46 = bb_auto_cover_out[691];
  assign coverage_47 = bb_auto_cover_out[690];
  assign coverage_48 = bb_auto_cover_out[689];
  assign coverage_49 = bb_auto_cover_out[688];
  assign coverage_50 = bb_auto_cover_out[687];
  assign coverage_51 = bb_auto_cover_out[686];
  assign coverage_52 = bb_auto_cover_out[332];
  assign coverage_53 = bb_auto_cover_out[331];
  assign coverage_54 = bb_auto_cover_out[330];
  assign coverage_55 = bb_auto_cover_out[329];
  assign coverage_56 = bb_auto_cover_out[328];
  assign coverage_57 = bb_auto_cover_out[327];
  assign coverage_58 = bb_auto_cover_out[326];
  assign coverage_59 = bb_auto_cover_out[325];
  assign coverage_60 = bb_auto_cover_out[324];
  assign coverage_61 = bb_auto_cover_out[323];
  assign coverage_62 = bb_auto_cover_out[322];
  assign coverage_63 = bb_auto_cover_out[321];
  assign coverage_64 = bb_auto_cover_out[320];
  assign coverage_65 = bb_auto_cover_out[319];
  assign coverage_66 = bb_auto_cover_out[318];
  assign coverage_67 = bb_auto_cover_out[317];
  assign coverage_68 = bb_auto_cover_out[316];
  assign coverage_69 = bb_auto_cover_out[309];
  assign coverage_70 = bb_auto_cover_out[304];
  assign coverage_71 = bb_auto_cover_out[303];
  assign coverage_72 = bb_auto_cover_out[302];
  assign coverage_73 = bb_auto_cover_out[301];
  assign coverage_74 = bb_auto_cover_out[300];
  assign coverage_75 = bb_auto_cover_out[299];
  assign coverage_76 = bb_auto_cover_out[298];
  assign coverage_77 = bb_auto_cover_out[297];
  assign coverage_78 = bb_auto_cover_out[295];
  assign coverage_79 = bb_auto_cover_out[294];
  assign coverage_80 = bb_auto_cover_out[291];
  assign coverage_81 = bb_auto_cover_out[290];
  assign coverage_82 = bb_auto_cover_out[289];
  assign coverage_83 = bb_auto_cover_out[285];
  assign coverage_84 = bb_auto_cover_out[281];
  assign coverage_85 = bb_auto_cover_out[279];
  assign coverage_86 = bb_auto_cover_out[278];
  assign coverage_87 = bb_auto_cover_out[277];
  assign coverage_88 = bb_auto_cover_out[276];
  assign coverage_89 = bb_auto_cover_out[275];
  assign coverage_90 = bb_auto_cover_out[274];
  assign coverage_91 = bb_auto_cover_out[273];
  assign coverage_92 = bb_auto_cover_out[272];
  assign coverage_93 = bb_auto_cover_out[271];
  assign coverage_94 = bb_auto_cover_out[270];
  assign coverage_95 = bb_auto_cover_out[269];
  assign coverage_96 = bb_auto_cover_out[268];
  assign coverage_97 = bb_auto_cover_out[267];
  assign coverage_98 = bb_auto_cover_out[266];
  assign coverage_99 = bb_auto_cover_out[265];
  assign coverage_100 = bb_auto_cover_out[264];
  assign coverage_101 = bb_auto_cover_out[263];
  assign coverage_102 = bb_auto_cover_out[262];
  assign coverage_103 = bb_auto_cover_out[261];
  assign coverage_104 = bb_auto_cover_out[260];
  assign coverage_105 = bb_auto_cover_out[259];
  assign coverage_106 = bb_auto_cover_out[258];
  assign coverage_107 = bb_auto_cover_out[257];
  assign coverage_108 = bb_auto_cover_out[256];
  assign coverage_109 = bb_auto_cover_out[255];
  assign coverage_110 = bb_auto_cover_out[254];
  assign coverage_111 = bb_auto_cover_out[253];
  assign coverage_112 = bb_auto_cover_out[252];
  assign coverage_113 = bb_auto_cover_out[251];
  assign coverage_114 = bb_auto_cover_out[250];
  assign coverage_115 = bb_auto_cover_out[249];
  assign coverage_116 = bb_auto_cover_out[248];
  assign coverage_117 = bb_auto_cover_out[247];
  assign coverage_118 = bb_auto_cover_out[246];
  assign coverage_119 = bb_auto_cover_out[245];
  assign coverage_120 = bb_auto_cover_out[244];
  assign coverage_121 = bb_auto_cover_out[243];
  assign coverage_122 = bb_auto_cover_out[242];
  assign coverage_123 = bb_auto_cover_out[241];
  assign coverage_124 = bb_auto_cover_out[240];
  assign coverage_125 = bb_auto_cover_out[239];
  assign coverage_126 = bb_auto_cover_out[238];
  assign coverage_127 = bb_auto_cover_out[237];
  assign coverage_128 = bb_auto_cover_out[236];
  assign coverage_129 = bb_auto_cover_out[235];
  assign coverage_130 = bb_auto_cover_out[234];
  assign coverage_131 = bb_auto_cover_out[233];
  assign coverage_132 = bb_auto_cover_out[232];
  assign coverage_133 = bb_auto_cover_out[231];
  assign coverage_134 = bb_auto_cover_out[230];
  assign coverage_135 = bb_auto_cover_out[229];
  assign coverage_136 = bb_auto_cover_out[228];
  assign coverage_137 = bb_auto_cover_out[227];
  assign coverage_138 = bb_auto_cover_out[226];
  assign coverage_139 = bb_auto_cover_out[225];
  assign coverage_140 = bb_auto_cover_out[224];
  assign coverage_141 = bb_auto_cover_out[223];
  assign coverage_142 = bb_auto_cover_out[222];
  assign coverage_143 = bb_auto_cover_out[221];
  assign coverage_144 = bb_auto_cover_out[220];
  assign coverage_145 = bb_auto_cover_out[219];
  assign coverage_146 = bb_auto_cover_out[218];
  assign coverage_147 = bb_auto_cover_out[217];
  assign coverage_148 = bb_auto_cover_out[216];
  assign coverage_149 = bb_auto_cover_out[215];
  assign coverage_150 = bb_auto_cover_out[214];
  assign coverage_151 = bb_auto_cover_out[213];
  assign coverage_152 = bb_auto_cover_out[212];
  assign coverage_153 = bb_auto_cover_out[211];
  assign coverage_154 = bb_auto_cover_out[210];
  assign coverage_155 = bb_auto_cover_out[209];
  assign coverage_156 = bb_auto_cover_out[208];
  assign coverage_157 = bb_auto_cover_out[207];
  assign coverage_158 = bb_auto_cover_out[206];
  assign coverage_159 = bb_auto_cover_out[205];
  assign coverage_160 = bb_auto_cover_out[204];
  assign coverage_161 = bb_auto_cover_out[203];
  assign coverage_162 = bb_auto_cover_out[202];
  assign coverage_163 = bb_auto_cover_out[201];
  assign coverage_164 = bb_auto_cover_out[200];
  assign coverage_165 = bb_auto_cover_out[199];
  assign coverage_166 = bb_auto_cover_out[198];
  assign coverage_167 = bb_auto_cover_out[126];
  assign coverage_168 = bb_auto_cover_out[122];
  assign coverage_169 = bb_auto_cover_out[111];
  assign coverage_170 = bb_auto_cover_out[47];
  assign coverage_171 = bb_auto_cover_out[46];
  assign coverage_172 = bb_auto_cover_out[45];
  assign coverage_173 = bb_auto_cover_out[44];
  assign coverage_174 = bb_auto_cover_out[43];
  assign coverage_175 = bb_auto_cover_out[42];
  assign coverage_176 = bb_auto_cover_out[41];
  assign coverage_177 = bb_auto_cover_out[40];
  assign coverage_178 = bb_auto_cover_out[39];
  assign coverage_179 = bb_auto_cover_out[38];
  assign coverage_180 = bb_auto_cover_out[37];
  assign coverage_181 = bb_auto_cover_out[36];
  assign coverage_182 = bb_auto_cover_out[34];
  assign coverage_183 = bb_auto_cover_out[33];
  assign coverage_184 = bb_auto_cover_out[32];
  assign coverage_185 = bb_auto_cover_out[31];
  assign coverage_186 = bb_auto_cover_out[24];
  assign coverage_187 = bb_auto_cover_out[23];
  assign coverage_188 = bb_auto_cover_out[19];
  assign coverage_189 = bb_auto_cover_out[7];
  assign coverage_190 = bb_auto_cover_out[6];
  assign coverage_191 = bb_auto_cover_out[2];
  assign io_coverage_0 = coverage_0;
  assign io_coverage_1 = coverage_1;
  assign io_coverage_2 = coverage_2;
  assign io_coverage_3 = coverage_3;
  assign io_coverage_4 = coverage_4;
  assign io_coverage_5 = coverage_5;
  assign io_coverage_6 = coverage_6;
  assign io_coverage_7 = coverage_7;
  assign io_coverage_8 = coverage_8;
  assign io_coverage_9 = coverage_9;
  assign io_coverage_10 = coverage_10;
  assign io_coverage_11 = coverage_11;
  assign io_coverage_12 = coverage_12;
  assign io_coverage_13 = coverage_13;
  assign io_coverage_14 = coverage_14;
  assign io_coverage_15 = coverage_15;
  assign io_coverage_16 = coverage_16;
  assign io_coverage_17 = coverage_17;
  assign io_coverage_18 = coverage_18;
  assign io_coverage_19 = coverage_19;
  assign io_coverage_20 = coverage_20;
  assign io_coverage_21 = coverage_21;
  assign io_coverage_22 = coverage_22;
  assign io_coverage_23 = coverage_23;
  assign io_coverage_24 = coverage_24;
  assign io_coverage_25 = coverage_25;
  assign io_coverage_26 = coverage_26;
  assign io_coverage_27 = coverage_27;
  assign io_coverage_28 = coverage_28;
  assign io_coverage_29 = coverage_29;
  assign io_coverage_30 = coverage_30;
  assign io_coverage_31 = coverage_31;
  assign io_coverage_32 = coverage_32;
  assign io_coverage_33 = coverage_33;
  assign io_coverage_34 = coverage_34;
  assign io_coverage_35 = coverage_35;
  assign io_coverage_36 = coverage_36;
  assign io_coverage_37 = coverage_37;
  assign io_coverage_38 = coverage_38;
  assign io_coverage_39 = coverage_39;
  assign io_coverage_40 = coverage_40;
  assign io_coverage_41 = coverage_41;
  assign io_coverage_42 = coverage_42;
  assign io_coverage_43 = coverage_43;
  assign io_coverage_44 = coverage_44;
  assign io_coverage_45 = coverage_45;
  assign io_coverage_46 = coverage_46;
  assign io_coverage_47 = coverage_47;
  assign io_coverage_48 = coverage_48;
  assign io_coverage_49 = coverage_49;
  assign io_coverage_50 = coverage_50;
  assign io_coverage_51 = coverage_51;
  assign io_coverage_52 = coverage_52;
  assign io_coverage_53 = coverage_53;
  assign io_coverage_54 = coverage_54;
  assign io_coverage_55 = coverage_55;
  assign io_coverage_56 = coverage_56;
  assign io_coverage_57 = coverage_57;
  assign io_coverage_58 = coverage_58;
  assign io_coverage_59 = coverage_59;
  assign io_coverage_60 = coverage_60;
  assign io_coverage_61 = coverage_61;
  assign io_coverage_62 = coverage_62;
  assign io_coverage_63 = coverage_63;
  assign io_coverage_64 = coverage_64;
  assign io_coverage_65 = coverage_65;
  assign io_coverage_66 = coverage_66;
  assign io_coverage_67 = coverage_67;
  assign io_coverage_68 = coverage_68;
  assign io_coverage_69 = coverage_69;
  assign io_coverage_70 = coverage_70;
  assign io_coverage_71 = coverage_71;
  assign io_coverage_72 = coverage_72;
  assign io_coverage_73 = coverage_73;
  assign io_coverage_74 = coverage_74;
  assign io_coverage_75 = coverage_75;
  assign io_coverage_76 = coverage_76;
  assign io_coverage_77 = coverage_77;
  assign io_coverage_78 = coverage_78;
  assign io_coverage_79 = coverage_79;
  assign io_coverage_80 = coverage_80;
  assign io_coverage_81 = coverage_81;
  assign io_coverage_82 = coverage_82;
  assign io_coverage_83 = coverage_83;
  assign io_coverage_84 = coverage_84;
  assign io_coverage_85 = coverage_85;
  assign io_coverage_86 = coverage_86;
  assign io_coverage_87 = coverage_87;
  assign io_coverage_88 = coverage_88;
  assign io_coverage_89 = coverage_89;
  assign io_coverage_90 = coverage_90;
  assign io_coverage_91 = coverage_91;
  assign io_coverage_92 = coverage_92;
  assign io_coverage_93 = coverage_93;
  assign io_coverage_94 = coverage_94;
  assign io_coverage_95 = coverage_95;
  assign io_coverage_96 = coverage_96;
  assign io_coverage_97 = coverage_97;
  assign io_coverage_98 = coverage_98;
  assign io_coverage_99 = coverage_99;
  assign io_coverage_100 = coverage_100;
  assign io_coverage_101 = coverage_101;
  assign io_coverage_102 = coverage_102;
  assign io_coverage_103 = coverage_103;
  assign io_coverage_104 = coverage_104;
  assign io_coverage_105 = coverage_105;
  assign io_coverage_106 = coverage_106;
  assign io_coverage_107 = coverage_107;
  assign io_coverage_108 = coverage_108;
  assign io_coverage_109 = coverage_109;
  assign io_coverage_110 = coverage_110;
  assign io_coverage_111 = coverage_111;
  assign io_coverage_112 = coverage_112;
  assign io_coverage_113 = coverage_113;
  assign io_coverage_114 = coverage_114;
  assign io_coverage_115 = coverage_115;
  assign io_coverage_116 = coverage_116;
  assign io_coverage_117 = coverage_117;
  assign io_coverage_118 = coverage_118;
  assign io_coverage_119 = coverage_119;
  assign io_coverage_120 = coverage_120;
  assign io_coverage_121 = coverage_121;
  assign io_coverage_122 = coverage_122;
  assign io_coverage_123 = coverage_123;
  assign io_coverage_124 = coverage_124;
  assign io_coverage_125 = coverage_125;
  assign io_coverage_126 = coverage_126;
  assign io_coverage_127 = coverage_127;
  assign io_coverage_128 = coverage_128;
  assign io_coverage_129 = coverage_129;
  assign io_coverage_130 = coverage_130;
  assign io_coverage_131 = coverage_131;
  assign io_coverage_132 = coverage_132;
  assign io_coverage_133 = coverage_133;
  assign io_coverage_134 = coverage_134;
  assign io_coverage_135 = coverage_135;
  assign io_coverage_136 = coverage_136;
  assign io_coverage_137 = coverage_137;
  assign io_coverage_138 = coverage_138;
  assign io_coverage_139 = coverage_139;
  assign io_coverage_140 = coverage_140;
  assign io_coverage_141 = coverage_141;
  assign io_coverage_142 = coverage_142;
  assign io_coverage_143 = coverage_143;
  assign io_coverage_144 = coverage_144;
  assign io_coverage_145 = coverage_145;
  assign io_coverage_146 = coverage_146;
  assign io_coverage_147 = coverage_147;
  assign io_coverage_148 = coverage_148;
  assign io_coverage_149 = coverage_149;
  assign io_coverage_150 = coverage_150;
  assign io_coverage_151 = coverage_151;
  assign io_coverage_152 = coverage_152;
  assign io_coverage_153 = coverage_153;
  assign io_coverage_154 = coverage_154;
  assign io_coverage_155 = coverage_155;
  assign io_coverage_156 = coverage_156;
  assign io_coverage_157 = coverage_157;
  assign io_coverage_158 = coverage_158;
  assign io_coverage_159 = coverage_159;
  assign io_coverage_160 = coverage_160;
  assign io_coverage_161 = coverage_161;
  assign io_coverage_162 = coverage_162;
  assign io_coverage_163 = coverage_163;
  assign io_coverage_164 = coverage_164;
  assign io_coverage_165 = coverage_165;
  assign io_coverage_166 = coverage_166;
  assign io_coverage_167 = coverage_167;
  assign io_coverage_168 = coverage_168;
  assign io_coverage_169 = coverage_169;
  assign io_coverage_170 = coverage_170;
  assign io_coverage_171 = coverage_171;
  assign io_coverage_172 = coverage_172;
  assign io_coverage_173 = coverage_173;
  assign io_coverage_174 = coverage_174;
  assign io_coverage_175 = coverage_175;
  assign io_coverage_176 = coverage_176;
  assign io_coverage_177 = coverage_177;
  assign io_coverage_178 = coverage_178;
  assign io_coverage_179 = coverage_179;
  assign io_coverage_180 = coverage_180;
  assign io_coverage_181 = coverage_181;
  assign io_coverage_182 = coverage_182;
  assign io_coverage_183 = coverage_183;
  assign io_coverage_184 = coverage_184;
  assign io_coverage_185 = coverage_185;
  assign io_coverage_186 = coverage_186;
  assign io_coverage_187 = coverage_187;
  assign io_coverage_188 = coverage_188;
  assign io_coverage_189 = coverage_189;
  assign io_coverage_190 = coverage_190;
  assign io_coverage_191 = coverage_191;
  assign bb_clock = clock;
  assign bb_reset = reset;
  assign bb_metaReset = io_meta_reset;
  assign bb_io_imem_resp_bits_data = _T_202;
  assign bb_io_imem_req_ready = _T_203;
  assign bb_io_imem_resp_valid = _T_204;
  assign bb_io_reset = _T_205;
endmodule
module SaturatingCounter(
  input   clock,
  input   reset,
  input   io_enable,
  output  io_value
);
  reg  count;
  reg [31:0] _RAND_0;
  wire  _T_7;
  wire  _T_9;
  wire [1:0] _T_11;
  wire  _T_12;
  wire  _T_13;
  assign _T_7 = io_enable == 1'h0;
  assign _T_9 = _T_7 | count;
  assign _T_11 = count + 1'h1;
  assign _T_12 = _T_11[0:0];
  assign _T_13 = _T_9 ? count : _T_12;
  assign io_value = count;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  count = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 1'h0;
    end else begin
      if (!(_T_9)) begin
        count <= _T_12;
      end
    end
  end
endmodule
module E2ECoverageHarness(
  input        clock,
  input        reset,
  input  [7:0] io_input_bytes_0,
  input  [7:0] io_input_bytes_1,
  input  [7:0] io_input_bytes_2,
  input  [7:0] io_input_bytes_3,
  input  [7:0] io_input_bytes_4,
  input  [7:0] io_input_bytes_5,
  input  [7:0] io_input_bytes_6,
  input  [7:0] io_input_bytes_7,
  output [7:0] io_coverage_bytes_0,
  output [7:0] io_coverage_bytes_1,
  output [7:0] io_coverage_bytes_2,
  output [7:0] io_coverage_bytes_3,
  output [7:0] io_coverage_bytes_4,
  output [7:0] io_coverage_bytes_5,
  output [7:0] io_coverage_bytes_6,
  output [7:0] io_coverage_bytes_7,
  output [7:0] io_coverage_bytes_8,
  output [7:0] io_coverage_bytes_9,
  output [7:0] io_coverage_bytes_10,
  output [7:0] io_coverage_bytes_11,
  output [7:0] io_coverage_bytes_12,
  output [7:0] io_coverage_bytes_13,
  output [7:0] io_coverage_bytes_14,
  output [7:0] io_coverage_bytes_15,
  output [7:0] io_coverage_bytes_16,
  output [7:0] io_coverage_bytes_17,
  output [7:0] io_coverage_bytes_18,
  output [7:0] io_coverage_bytes_19,
  output [7:0] io_coverage_bytes_20,
  output [7:0] io_coverage_bytes_21,
  output [7:0] io_coverage_bytes_22,
  output [7:0] io_coverage_bytes_23,
  output [7:0] io_coverage_bytes_24,
  output [7:0] io_coverage_bytes_25,
  output [7:0] io_coverage_bytes_26,
  output [7:0] io_coverage_bytes_27,
  output [7:0] io_coverage_bytes_28,
  output [7:0] io_coverage_bytes_29,
  output [7:0] io_coverage_bytes_30,
  output [7:0] io_coverage_bytes_31,
  output [7:0] io_coverage_bytes_32,
  output [7:0] io_coverage_bytes_33,
  output [7:0] io_coverage_bytes_34,
  output [7:0] io_coverage_bytes_35,
  output [7:0] io_coverage_bytes_36,
  output [7:0] io_coverage_bytes_37,
  output [7:0] io_coverage_bytes_38,
  output [7:0] io_coverage_bytes_39,
  output [7:0] io_coverage_bytes_40,
  output [7:0] io_coverage_bytes_41,
  output [7:0] io_coverage_bytes_42,
  output [7:0] io_coverage_bytes_43,
  output [7:0] io_coverage_bytes_44,
  output [7:0] io_coverage_bytes_45,
  output [7:0] io_coverage_bytes_46,
  output [7:0] io_coverage_bytes_47,
  output [7:0] io_coverage_bytes_48,
  output [7:0] io_coverage_bytes_49,
  output [7:0] io_coverage_bytes_50,
  output [7:0] io_coverage_bytes_51,
  output [7:0] io_coverage_bytes_52,
  output [7:0] io_coverage_bytes_53,
  output [7:0] io_coverage_bytes_54,
  output [7:0] io_coverage_bytes_55,
  output [7:0] io_coverage_bytes_56,
  output [7:0] io_coverage_bytes_57,
  output [7:0] io_coverage_bytes_58,
  output [7:0] io_coverage_bytes_59,
  output [7:0] io_coverage_bytes_60,
  output [7:0] io_coverage_bytes_61,
  output [7:0] io_coverage_bytes_62,
  output [7:0] io_coverage_bytes_63,
  output [7:0] io_coverage_bytes_64,
  output [7:0] io_coverage_bytes_65,
  output [7:0] io_coverage_bytes_66,
  output [7:0] io_coverage_bytes_67,
  output [7:0] io_coverage_bytes_68,
  output [7:0] io_coverage_bytes_69,
  output [7:0] io_coverage_bytes_70,
  output [7:0] io_coverage_bytes_71,
  output [7:0] io_coverage_bytes_72,
  output [7:0] io_coverage_bytes_73,
  output [7:0] io_coverage_bytes_74,
  output [7:0] io_coverage_bytes_75,
  output [7:0] io_coverage_bytes_76,
  output [7:0] io_coverage_bytes_77,
  output [7:0] io_coverage_bytes_78,
  output [7:0] io_coverage_bytes_79,
  output [7:0] io_coverage_bytes_80,
  output [7:0] io_coverage_bytes_81,
  output [7:0] io_coverage_bytes_82,
  output [7:0] io_coverage_bytes_83,
  output [7:0] io_coverage_bytes_84,
  output [7:0] io_coverage_bytes_85,
  output [7:0] io_coverage_bytes_86,
  output [7:0] io_coverage_bytes_87,
  output [7:0] io_coverage_bytes_88,
  output [7:0] io_coverage_bytes_89,
  output [7:0] io_coverage_bytes_90,
  output [7:0] io_coverage_bytes_91,
  output [7:0] io_coverage_bytes_92,
  output [7:0] io_coverage_bytes_93,
  output [7:0] io_coverage_bytes_94,
  output [7:0] io_coverage_bytes_95,
  output [7:0] io_coverage_bytes_96,
  output [7:0] io_coverage_bytes_97,
  output [7:0] io_coverage_bytes_98,
  output [7:0] io_coverage_bytes_99,
  output [7:0] io_coverage_bytes_100,
  output [7:0] io_coverage_bytes_101,
  output [7:0] io_coverage_bytes_102,
  output [7:0] io_coverage_bytes_103,
  output [7:0] io_coverage_bytes_104,
  output [7:0] io_coverage_bytes_105,
  output [7:0] io_coverage_bytes_106,
  output [7:0] io_coverage_bytes_107,
  output [7:0] io_coverage_bytes_108,
  output [7:0] io_coverage_bytes_109,
  output [7:0] io_coverage_bytes_110,
  output [7:0] io_coverage_bytes_111,
  output [7:0] io_coverage_bytes_112,
  output [7:0] io_coverage_bytes_113,
  output [7:0] io_coverage_bytes_114,
  output [7:0] io_coverage_bytes_115,
  output [7:0] io_coverage_bytes_116,
  output [7:0] io_coverage_bytes_117,
  output [7:0] io_coverage_bytes_118,
  output [7:0] io_coverage_bytes_119,
  output [7:0] io_coverage_bytes_120,
  output [7:0] io_coverage_bytes_121,
  output [7:0] io_coverage_bytes_122,
  output [7:0] io_coverage_bytes_123,
  output [7:0] io_coverage_bytes_124,
  output [7:0] io_coverage_bytes_125,
  output [7:0] io_coverage_bytes_126,
  output [7:0] io_coverage_bytes_127,
  output [7:0] io_coverage_bytes_128,
  output [7:0] io_coverage_bytes_129,
  output [7:0] io_coverage_bytes_130,
  output [7:0] io_coverage_bytes_131,
  output [7:0] io_coverage_bytes_132,
  output [7:0] io_coverage_bytes_133,
  output [7:0] io_coverage_bytes_134,
  output [7:0] io_coverage_bytes_135,
  output [7:0] io_coverage_bytes_136,
  output [7:0] io_coverage_bytes_137,
  output [7:0] io_coverage_bytes_138,
  output [7:0] io_coverage_bytes_139,
  output [7:0] io_coverage_bytes_140,
  output [7:0] io_coverage_bytes_141,
  output [7:0] io_coverage_bytes_142,
  output [7:0] io_coverage_bytes_143,
  output [7:0] io_coverage_bytes_144,
  output [7:0] io_coverage_bytes_145,
  output [7:0] io_coverage_bytes_146,
  output [7:0] io_coverage_bytes_147,
  output [7:0] io_coverage_bytes_148,
  output [7:0] io_coverage_bytes_149,
  output [7:0] io_coverage_bytes_150,
  output [7:0] io_coverage_bytes_151,
  output [7:0] io_coverage_bytes_152,
  output [7:0] io_coverage_bytes_153,
  output [7:0] io_coverage_bytes_154,
  output [7:0] io_coverage_bytes_155,
  output [7:0] io_coverage_bytes_156,
  output [7:0] io_coverage_bytes_157,
  output [7:0] io_coverage_bytes_158,
  output [7:0] io_coverage_bytes_159,
  output [7:0] io_coverage_bytes_160,
  output [7:0] io_coverage_bytes_161,
  output [7:0] io_coverage_bytes_162,
  output [7:0] io_coverage_bytes_163,
  output [7:0] io_coverage_bytes_164,
  output [7:0] io_coverage_bytes_165,
  output [7:0] io_coverage_bytes_166,
  output [7:0] io_coverage_bytes_167,
  output [7:0] io_coverage_bytes_168,
  output [7:0] io_coverage_bytes_169,
  output [7:0] io_coverage_bytes_170,
  output [7:0] io_coverage_bytes_171,
  output [7:0] io_coverage_bytes_172,
  output [7:0] io_coverage_bytes_173,
  output [7:0] io_coverage_bytes_174,
  output [7:0] io_coverage_bytes_175,
  output [7:0] io_coverage_bytes_176,
  output [7:0] io_coverage_bytes_177,
  output [7:0] io_coverage_bytes_178,
  output [7:0] io_coverage_bytes_179,
  output [7:0] io_coverage_bytes_180,
  output [7:0] io_coverage_bytes_181,
  output [7:0] io_coverage_bytes_182,
  output [7:0] io_coverage_bytes_183,
  output [7:0] io_coverage_bytes_184,
  output [7:0] io_coverage_bytes_185,
  output [7:0] io_coverage_bytes_186,
  output [7:0] io_coverage_bytes_187,
  output [7:0] io_coverage_bytes_188,
  output [7:0] io_coverage_bytes_189,
  output [7:0] io_coverage_bytes_190,
  output [7:0] io_coverage_bytes_191,
  output [7:0] io_coverage_bytes_192,
  output [7:0] io_coverage_bytes_193,
  output [7:0] io_coverage_bytes_194,
  output [7:0] io_coverage_bytes_195,
  output [7:0] io_coverage_bytes_196,
  output [7:0] io_coverage_bytes_197,
  input        io_meta_reset
);
  wire  dut_clock;
  wire  dut_reset;
  wire  dut_io_meta_reset;
  wire [34:0] dut_io_inputs;
  wire  dut_io_coverage_0;
  wire  dut_io_coverage_1;
  wire  dut_io_coverage_2;
  wire  dut_io_coverage_3;
  wire  dut_io_coverage_4;
  wire  dut_io_coverage_5;
  wire  dut_io_coverage_6;
  wire  dut_io_coverage_7;
  wire  dut_io_coverage_8;
  wire  dut_io_coverage_9;
  wire  dut_io_coverage_10;
  wire  dut_io_coverage_11;
  wire  dut_io_coverage_12;
  wire  dut_io_coverage_13;
  wire  dut_io_coverage_14;
  wire  dut_io_coverage_15;
  wire  dut_io_coverage_16;
  wire  dut_io_coverage_17;
  wire  dut_io_coverage_18;
  wire  dut_io_coverage_19;
  wire  dut_io_coverage_20;
  wire  dut_io_coverage_21;
  wire  dut_io_coverage_22;
  wire  dut_io_coverage_23;
  wire  dut_io_coverage_24;
  wire  dut_io_coverage_25;
  wire  dut_io_coverage_26;
  wire  dut_io_coverage_27;
  wire  dut_io_coverage_28;
  wire  dut_io_coverage_29;
  wire  dut_io_coverage_30;
  wire  dut_io_coverage_31;
  wire  dut_io_coverage_32;
  wire  dut_io_coverage_33;
  wire  dut_io_coverage_34;
  wire  dut_io_coverage_35;
  wire  dut_io_coverage_36;
  wire  dut_io_coverage_37;
  wire  dut_io_coverage_38;
  wire  dut_io_coverage_39;
  wire  dut_io_coverage_40;
  wire  dut_io_coverage_41;
  wire  dut_io_coverage_42;
  wire  dut_io_coverage_43;
  wire  dut_io_coverage_44;
  wire  dut_io_coverage_45;
  wire  dut_io_coverage_46;
  wire  dut_io_coverage_47;
  wire  dut_io_coverage_48;
  wire  dut_io_coverage_49;
  wire  dut_io_coverage_50;
  wire  dut_io_coverage_51;
  wire  dut_io_coverage_52;
  wire  dut_io_coverage_53;
  wire  dut_io_coverage_54;
  wire  dut_io_coverage_55;
  wire  dut_io_coverage_56;
  wire  dut_io_coverage_57;
  wire  dut_io_coverage_58;
  wire  dut_io_coverage_59;
  wire  dut_io_coverage_60;
  wire  dut_io_coverage_61;
  wire  dut_io_coverage_62;
  wire  dut_io_coverage_63;
  wire  dut_io_coverage_64;
  wire  dut_io_coverage_65;
  wire  dut_io_coverage_66;
  wire  dut_io_coverage_67;
  wire  dut_io_coverage_68;
  wire  dut_io_coverage_69;
  wire  dut_io_coverage_70;
  wire  dut_io_coverage_71;
  wire  dut_io_coverage_72;
  wire  dut_io_coverage_73;
  wire  dut_io_coverage_74;
  wire  dut_io_coverage_75;
  wire  dut_io_coverage_76;
  wire  dut_io_coverage_77;
  wire  dut_io_coverage_78;
  wire  dut_io_coverage_79;
  wire  dut_io_coverage_80;
  wire  dut_io_coverage_81;
  wire  dut_io_coverage_82;
  wire  dut_io_coverage_83;
  wire  dut_io_coverage_84;
  wire  dut_io_coverage_85;
  wire  dut_io_coverage_86;
  wire  dut_io_coverage_87;
  wire  dut_io_coverage_88;
  wire  dut_io_coverage_89;
  wire  dut_io_coverage_90;
  wire  dut_io_coverage_91;
  wire  dut_io_coverage_92;
  wire  dut_io_coverage_93;
  wire  dut_io_coverage_94;
  wire  dut_io_coverage_95;
  wire  dut_io_coverage_96;
  wire  dut_io_coverage_97;
  wire  dut_io_coverage_98;
  wire  dut_io_coverage_99;
  wire  dut_io_coverage_100;
  wire  dut_io_coverage_101;
  wire  dut_io_coverage_102;
  wire  dut_io_coverage_103;
  wire  dut_io_coverage_104;
  wire  dut_io_coverage_105;
  wire  dut_io_coverage_106;
  wire  dut_io_coverage_107;
  wire  dut_io_coverage_108;
  wire  dut_io_coverage_109;
  wire  dut_io_coverage_110;
  wire  dut_io_coverage_111;
  wire  dut_io_coverage_112;
  wire  dut_io_coverage_113;
  wire  dut_io_coverage_114;
  wire  dut_io_coverage_115;
  wire  dut_io_coverage_116;
  wire  dut_io_coverage_117;
  wire  dut_io_coverage_118;
  wire  dut_io_coverage_119;
  wire  dut_io_coverage_120;
  wire  dut_io_coverage_121;
  wire  dut_io_coverage_122;
  wire  dut_io_coverage_123;
  wire  dut_io_coverage_124;
  wire  dut_io_coverage_125;
  wire  dut_io_coverage_126;
  wire  dut_io_coverage_127;
  wire  dut_io_coverage_128;
  wire  dut_io_coverage_129;
  wire  dut_io_coverage_130;
  wire  dut_io_coverage_131;
  wire  dut_io_coverage_132;
  wire  dut_io_coverage_133;
  wire  dut_io_coverage_134;
  wire  dut_io_coverage_135;
  wire  dut_io_coverage_136;
  wire  dut_io_coverage_137;
  wire  dut_io_coverage_138;
  wire  dut_io_coverage_139;
  wire  dut_io_coverage_140;
  wire  dut_io_coverage_141;
  wire  dut_io_coverage_142;
  wire  dut_io_coverage_143;
  wire  dut_io_coverage_144;
  wire  dut_io_coverage_145;
  wire  dut_io_coverage_146;
  wire  dut_io_coverage_147;
  wire  dut_io_coverage_148;
  wire  dut_io_coverage_149;
  wire  dut_io_coverage_150;
  wire  dut_io_coverage_151;
  wire  dut_io_coverage_152;
  wire  dut_io_coverage_153;
  wire  dut_io_coverage_154;
  wire  dut_io_coverage_155;
  wire  dut_io_coverage_156;
  wire  dut_io_coverage_157;
  wire  dut_io_coverage_158;
  wire  dut_io_coverage_159;
  wire  dut_io_coverage_160;
  wire  dut_io_coverage_161;
  wire  dut_io_coverage_162;
  wire  dut_io_coverage_163;
  wire  dut_io_coverage_164;
  wire  dut_io_coverage_165;
  wire  dut_io_coverage_166;
  wire  dut_io_coverage_167;
  wire  dut_io_coverage_168;
  wire  dut_io_coverage_169;
  wire  dut_io_coverage_170;
  wire  dut_io_coverage_171;
  wire  dut_io_coverage_172;
  wire  dut_io_coverage_173;
  wire  dut_io_coverage_174;
  wire  dut_io_coverage_175;
  wire  dut_io_coverage_176;
  wire  dut_io_coverage_177;
  wire  dut_io_coverage_178;
  wire  dut_io_coverage_179;
  wire  dut_io_coverage_180;
  wire  dut_io_coverage_181;
  wire  dut_io_coverage_182;
  wire  dut_io_coverage_183;
  wire  dut_io_coverage_184;
  wire  dut_io_coverage_185;
  wire  dut_io_coverage_186;
  wire  dut_io_coverage_187;
  wire  dut_io_coverage_188;
  wire  dut_io_coverage_189;
  wire  dut_io_coverage_190;
  wire  dut_io_coverage_191;
  wire [15:0] _T_219;
  wire [15:0] _T_220;
  wire [31:0] _T_221;
  wire [15:0] _T_222;
  wire [15:0] _T_223;
  wire [31:0] _T_224;
  wire [63:0] input_bytes;
  wire [34:0] _T_225;
  wire  _T_227;
  wire  SaturatingCounter_clock;
  wire  SaturatingCounter_reset;
  wire  SaturatingCounter_io_enable;
  wire  SaturatingCounter_io_value;
  wire [7:0] coverage_0;
  wire  SaturatingCounter_1_clock;
  wire  SaturatingCounter_1_reset;
  wire  SaturatingCounter_1_io_enable;
  wire  SaturatingCounter_1_io_value;
  wire  _T_232;
  wire  SaturatingCounter_2_clock;
  wire  SaturatingCounter_2_reset;
  wire  SaturatingCounter_2_io_enable;
  wire  SaturatingCounter_2_io_value;
  wire  _T_233;
  wire [6:0] _T_237;
  wire [7:0] coverage_1;
  wire  SaturatingCounter_3_clock;
  wire  SaturatingCounter_3_reset;
  wire  SaturatingCounter_3_io_enable;
  wire  SaturatingCounter_3_io_value;
  wire  _T_239;
  wire  SaturatingCounter_4_clock;
  wire  SaturatingCounter_4_reset;
  wire  SaturatingCounter_4_io_enable;
  wire  SaturatingCounter_4_io_value;
  wire  _T_240;
  wire [6:0] _T_244;
  wire [7:0] coverage_2;
  wire  SaturatingCounter_5_clock;
  wire  SaturatingCounter_5_reset;
  wire  SaturatingCounter_5_io_enable;
  wire  SaturatingCounter_5_io_value;
  wire  _T_246;
  wire  SaturatingCounter_6_clock;
  wire  SaturatingCounter_6_reset;
  wire  SaturatingCounter_6_io_enable;
  wire  SaturatingCounter_6_io_value;
  wire  _T_247;
  wire [6:0] _T_251;
  wire [7:0] coverage_3;
  wire  SaturatingCounter_7_clock;
  wire  SaturatingCounter_7_reset;
  wire  SaturatingCounter_7_io_enable;
  wire  SaturatingCounter_7_io_value;
  wire  _T_253;
  wire  SaturatingCounter_8_clock;
  wire  SaturatingCounter_8_reset;
  wire  SaturatingCounter_8_io_enable;
  wire  SaturatingCounter_8_io_value;
  wire  _T_254;
  wire [6:0] _T_258;
  wire [7:0] coverage_4;
  wire  SaturatingCounter_9_clock;
  wire  SaturatingCounter_9_reset;
  wire  SaturatingCounter_9_io_enable;
  wire  SaturatingCounter_9_io_value;
  wire  _T_260;
  wire  SaturatingCounter_10_clock;
  wire  SaturatingCounter_10_reset;
  wire  SaturatingCounter_10_io_enable;
  wire  SaturatingCounter_10_io_value;
  wire  _T_261;
  wire [6:0] _T_265;
  wire [7:0] coverage_5;
  wire  SaturatingCounter_11_clock;
  wire  SaturatingCounter_11_reset;
  wire  SaturatingCounter_11_io_enable;
  wire  SaturatingCounter_11_io_value;
  wire  _T_267;
  wire  SaturatingCounter_12_clock;
  wire  SaturatingCounter_12_reset;
  wire  SaturatingCounter_12_io_enable;
  wire  SaturatingCounter_12_io_value;
  wire  _T_268;
  wire [6:0] _T_272;
  wire [7:0] coverage_6;
  wire  SaturatingCounter_13_clock;
  wire  SaturatingCounter_13_reset;
  wire  SaturatingCounter_13_io_enable;
  wire  SaturatingCounter_13_io_value;
  wire  _T_274;
  wire  SaturatingCounter_14_clock;
  wire  SaturatingCounter_14_reset;
  wire  SaturatingCounter_14_io_enable;
  wire  SaturatingCounter_14_io_value;
  wire  _T_275;
  wire [6:0] _T_279;
  wire [7:0] coverage_7;
  wire  SaturatingCounter_15_clock;
  wire  SaturatingCounter_15_reset;
  wire  SaturatingCounter_15_io_enable;
  wire  SaturatingCounter_15_io_value;
  wire  _T_281;
  wire  SaturatingCounter_16_clock;
  wire  SaturatingCounter_16_reset;
  wire  SaturatingCounter_16_io_enable;
  wire  SaturatingCounter_16_io_value;
  wire  _T_282;
  wire [6:0] _T_286;
  wire [7:0] coverage_8;
  wire  SaturatingCounter_17_clock;
  wire  SaturatingCounter_17_reset;
  wire  SaturatingCounter_17_io_enable;
  wire  SaturatingCounter_17_io_value;
  wire  _T_288;
  wire  SaturatingCounter_18_clock;
  wire  SaturatingCounter_18_reset;
  wire  SaturatingCounter_18_io_enable;
  wire  SaturatingCounter_18_io_value;
  wire  _T_289;
  wire [6:0] _T_293;
  wire [7:0] coverage_9;
  wire  SaturatingCounter_19_clock;
  wire  SaturatingCounter_19_reset;
  wire  SaturatingCounter_19_io_enable;
  wire  SaturatingCounter_19_io_value;
  wire  _T_295;
  wire  SaturatingCounter_20_clock;
  wire  SaturatingCounter_20_reset;
  wire  SaturatingCounter_20_io_enable;
  wire  SaturatingCounter_20_io_value;
  wire  _T_296;
  wire [6:0] _T_300;
  wire [7:0] coverage_10;
  wire  SaturatingCounter_21_clock;
  wire  SaturatingCounter_21_reset;
  wire  SaturatingCounter_21_io_enable;
  wire  SaturatingCounter_21_io_value;
  wire  _T_302;
  wire  SaturatingCounter_22_clock;
  wire  SaturatingCounter_22_reset;
  wire  SaturatingCounter_22_io_enable;
  wire  SaturatingCounter_22_io_value;
  wire  _T_303;
  wire [6:0] _T_307;
  wire [7:0] coverage_11;
  wire  SaturatingCounter_23_clock;
  wire  SaturatingCounter_23_reset;
  wire  SaturatingCounter_23_io_enable;
  wire  SaturatingCounter_23_io_value;
  wire  _T_309;
  wire  SaturatingCounter_24_clock;
  wire  SaturatingCounter_24_reset;
  wire  SaturatingCounter_24_io_enable;
  wire  SaturatingCounter_24_io_value;
  wire  _T_310;
  wire [6:0] _T_314;
  wire [7:0] coverage_12;
  wire  SaturatingCounter_25_clock;
  wire  SaturatingCounter_25_reset;
  wire  SaturatingCounter_25_io_enable;
  wire  SaturatingCounter_25_io_value;
  wire  _T_316;
  wire  SaturatingCounter_26_clock;
  wire  SaturatingCounter_26_reset;
  wire  SaturatingCounter_26_io_enable;
  wire  SaturatingCounter_26_io_value;
  wire  _T_317;
  wire [6:0] _T_321;
  wire [7:0] coverage_13;
  wire  SaturatingCounter_27_clock;
  wire  SaturatingCounter_27_reset;
  wire  SaturatingCounter_27_io_enable;
  wire  SaturatingCounter_27_io_value;
  wire  _T_323;
  wire  SaturatingCounter_28_clock;
  wire  SaturatingCounter_28_reset;
  wire  SaturatingCounter_28_io_enable;
  wire  SaturatingCounter_28_io_value;
  wire  _T_324;
  wire [6:0] _T_328;
  wire [7:0] coverage_14;
  wire  SaturatingCounter_29_clock;
  wire  SaturatingCounter_29_reset;
  wire  SaturatingCounter_29_io_enable;
  wire  SaturatingCounter_29_io_value;
  wire  _T_330;
  wire  SaturatingCounter_30_clock;
  wire  SaturatingCounter_30_reset;
  wire  SaturatingCounter_30_io_enable;
  wire  SaturatingCounter_30_io_value;
  wire  _T_331;
  wire [6:0] _T_335;
  wire [7:0] coverage_15;
  wire  SaturatingCounter_31_clock;
  wire  SaturatingCounter_31_reset;
  wire  SaturatingCounter_31_io_enable;
  wire  SaturatingCounter_31_io_value;
  wire  _T_337;
  wire  SaturatingCounter_32_clock;
  wire  SaturatingCounter_32_reset;
  wire  SaturatingCounter_32_io_enable;
  wire  SaturatingCounter_32_io_value;
  wire  _T_338;
  wire [6:0] _T_342;
  wire [7:0] coverage_16;
  wire  SaturatingCounter_33_clock;
  wire  SaturatingCounter_33_reset;
  wire  SaturatingCounter_33_io_enable;
  wire  SaturatingCounter_33_io_value;
  wire  _T_344;
  wire  SaturatingCounter_34_clock;
  wire  SaturatingCounter_34_reset;
  wire  SaturatingCounter_34_io_enable;
  wire  SaturatingCounter_34_io_value;
  wire  _T_345;
  wire [6:0] _T_349;
  wire [7:0] coverage_17;
  wire  SaturatingCounter_35_clock;
  wire  SaturatingCounter_35_reset;
  wire  SaturatingCounter_35_io_enable;
  wire  SaturatingCounter_35_io_value;
  wire  _T_351;
  wire  SaturatingCounter_36_clock;
  wire  SaturatingCounter_36_reset;
  wire  SaturatingCounter_36_io_enable;
  wire  SaturatingCounter_36_io_value;
  wire  _T_352;
  wire [6:0] _T_356;
  wire [7:0] coverage_18;
  wire  SaturatingCounter_37_clock;
  wire  SaturatingCounter_37_reset;
  wire  SaturatingCounter_37_io_enable;
  wire  SaturatingCounter_37_io_value;
  wire  _T_358;
  wire  SaturatingCounter_38_clock;
  wire  SaturatingCounter_38_reset;
  wire  SaturatingCounter_38_io_enable;
  wire  SaturatingCounter_38_io_value;
  wire  _T_359;
  wire [6:0] _T_363;
  wire [7:0] coverage_19;
  wire  SaturatingCounter_39_clock;
  wire  SaturatingCounter_39_reset;
  wire  SaturatingCounter_39_io_enable;
  wire  SaturatingCounter_39_io_value;
  wire  _T_365;
  wire  SaturatingCounter_40_clock;
  wire  SaturatingCounter_40_reset;
  wire  SaturatingCounter_40_io_enable;
  wire  SaturatingCounter_40_io_value;
  wire  _T_366;
  wire [6:0] _T_370;
  wire [7:0] coverage_20;
  wire  SaturatingCounter_41_clock;
  wire  SaturatingCounter_41_reset;
  wire  SaturatingCounter_41_io_enable;
  wire  SaturatingCounter_41_io_value;
  wire  _T_372;
  wire  SaturatingCounter_42_clock;
  wire  SaturatingCounter_42_reset;
  wire  SaturatingCounter_42_io_enable;
  wire  SaturatingCounter_42_io_value;
  wire  _T_373;
  wire [6:0] _T_377;
  wire [7:0] coverage_21;
  wire  SaturatingCounter_43_clock;
  wire  SaturatingCounter_43_reset;
  wire  SaturatingCounter_43_io_enable;
  wire  SaturatingCounter_43_io_value;
  wire  _T_379;
  wire  SaturatingCounter_44_clock;
  wire  SaturatingCounter_44_reset;
  wire  SaturatingCounter_44_io_enable;
  wire  SaturatingCounter_44_io_value;
  wire  _T_380;
  wire [6:0] _T_384;
  wire [7:0] coverage_22;
  wire  SaturatingCounter_45_clock;
  wire  SaturatingCounter_45_reset;
  wire  SaturatingCounter_45_io_enable;
  wire  SaturatingCounter_45_io_value;
  wire  _T_386;
  wire  SaturatingCounter_46_clock;
  wire  SaturatingCounter_46_reset;
  wire  SaturatingCounter_46_io_enable;
  wire  SaturatingCounter_46_io_value;
  wire  _T_387;
  wire [6:0] _T_391;
  wire [7:0] coverage_23;
  wire  SaturatingCounter_47_clock;
  wire  SaturatingCounter_47_reset;
  wire  SaturatingCounter_47_io_enable;
  wire  SaturatingCounter_47_io_value;
  wire  _T_393;
  wire  SaturatingCounter_48_clock;
  wire  SaturatingCounter_48_reset;
  wire  SaturatingCounter_48_io_enable;
  wire  SaturatingCounter_48_io_value;
  wire  _T_394;
  wire [6:0] _T_398;
  wire [7:0] coverage_24;
  wire  SaturatingCounter_49_clock;
  wire  SaturatingCounter_49_reset;
  wire  SaturatingCounter_49_io_enable;
  wire  SaturatingCounter_49_io_value;
  wire  _T_400;
  wire  SaturatingCounter_50_clock;
  wire  SaturatingCounter_50_reset;
  wire  SaturatingCounter_50_io_enable;
  wire  SaturatingCounter_50_io_value;
  wire  _T_401;
  wire [6:0] _T_405;
  wire [7:0] coverage_25;
  wire  SaturatingCounter_51_clock;
  wire  SaturatingCounter_51_reset;
  wire  SaturatingCounter_51_io_enable;
  wire  SaturatingCounter_51_io_value;
  wire  _T_407;
  wire  SaturatingCounter_52_clock;
  wire  SaturatingCounter_52_reset;
  wire  SaturatingCounter_52_io_enable;
  wire  SaturatingCounter_52_io_value;
  wire  _T_408;
  wire [6:0] _T_412;
  wire [7:0] coverage_26;
  wire  SaturatingCounter_53_clock;
  wire  SaturatingCounter_53_reset;
  wire  SaturatingCounter_53_io_enable;
  wire  SaturatingCounter_53_io_value;
  wire  _T_414;
  wire  SaturatingCounter_54_clock;
  wire  SaturatingCounter_54_reset;
  wire  SaturatingCounter_54_io_enable;
  wire  SaturatingCounter_54_io_value;
  wire  _T_415;
  wire [6:0] _T_419;
  wire [7:0] coverage_27;
  wire  SaturatingCounter_55_clock;
  wire  SaturatingCounter_55_reset;
  wire  SaturatingCounter_55_io_enable;
  wire  SaturatingCounter_55_io_value;
  wire  _T_421;
  wire  SaturatingCounter_56_clock;
  wire  SaturatingCounter_56_reset;
  wire  SaturatingCounter_56_io_enable;
  wire  SaturatingCounter_56_io_value;
  wire  _T_422;
  wire [6:0] _T_426;
  wire [7:0] coverage_28;
  wire  SaturatingCounter_57_clock;
  wire  SaturatingCounter_57_reset;
  wire  SaturatingCounter_57_io_enable;
  wire  SaturatingCounter_57_io_value;
  wire  _T_428;
  wire  SaturatingCounter_58_clock;
  wire  SaturatingCounter_58_reset;
  wire  SaturatingCounter_58_io_enable;
  wire  SaturatingCounter_58_io_value;
  wire  _T_429;
  wire [6:0] _T_433;
  wire [7:0] coverage_29;
  wire  SaturatingCounter_59_clock;
  wire  SaturatingCounter_59_reset;
  wire  SaturatingCounter_59_io_enable;
  wire  SaturatingCounter_59_io_value;
  wire  _T_435;
  wire  SaturatingCounter_60_clock;
  wire  SaturatingCounter_60_reset;
  wire  SaturatingCounter_60_io_enable;
  wire  SaturatingCounter_60_io_value;
  wire  _T_436;
  wire [6:0] _T_440;
  wire [7:0] coverage_30;
  wire  SaturatingCounter_61_clock;
  wire  SaturatingCounter_61_reset;
  wire  SaturatingCounter_61_io_enable;
  wire  SaturatingCounter_61_io_value;
  wire  _T_442;
  wire  SaturatingCounter_62_clock;
  wire  SaturatingCounter_62_reset;
  wire  SaturatingCounter_62_io_enable;
  wire  SaturatingCounter_62_io_value;
  wire  _T_443;
  wire [6:0] _T_447;
  wire [7:0] coverage_31;
  wire  SaturatingCounter_63_clock;
  wire  SaturatingCounter_63_reset;
  wire  SaturatingCounter_63_io_enable;
  wire  SaturatingCounter_63_io_value;
  wire  _T_449;
  wire  SaturatingCounter_64_clock;
  wire  SaturatingCounter_64_reset;
  wire  SaturatingCounter_64_io_enable;
  wire  SaturatingCounter_64_io_value;
  wire  _T_450;
  wire [6:0] _T_454;
  wire [7:0] coverage_32;
  wire  SaturatingCounter_65_clock;
  wire  SaturatingCounter_65_reset;
  wire  SaturatingCounter_65_io_enable;
  wire  SaturatingCounter_65_io_value;
  wire  _T_456;
  wire  SaturatingCounter_66_clock;
  wire  SaturatingCounter_66_reset;
  wire  SaturatingCounter_66_io_enable;
  wire  SaturatingCounter_66_io_value;
  wire  _T_457;
  wire [6:0] _T_461;
  wire [7:0] coverage_33;
  wire  SaturatingCounter_67_clock;
  wire  SaturatingCounter_67_reset;
  wire  SaturatingCounter_67_io_enable;
  wire  SaturatingCounter_67_io_value;
  wire  _T_463;
  wire  SaturatingCounter_68_clock;
  wire  SaturatingCounter_68_reset;
  wire  SaturatingCounter_68_io_enable;
  wire  SaturatingCounter_68_io_value;
  wire  _T_464;
  wire [6:0] _T_468;
  wire [7:0] coverage_34;
  wire  SaturatingCounter_69_clock;
  wire  SaturatingCounter_69_reset;
  wire  SaturatingCounter_69_io_enable;
  wire  SaturatingCounter_69_io_value;
  wire  _T_470;
  wire  SaturatingCounter_70_clock;
  wire  SaturatingCounter_70_reset;
  wire  SaturatingCounter_70_io_enable;
  wire  SaturatingCounter_70_io_value;
  wire  _T_471;
  wire [6:0] _T_475;
  wire [7:0] coverage_35;
  wire  SaturatingCounter_71_clock;
  wire  SaturatingCounter_71_reset;
  wire  SaturatingCounter_71_io_enable;
  wire  SaturatingCounter_71_io_value;
  wire  _T_477;
  wire  SaturatingCounter_72_clock;
  wire  SaturatingCounter_72_reset;
  wire  SaturatingCounter_72_io_enable;
  wire  SaturatingCounter_72_io_value;
  wire  _T_478;
  wire [6:0] _T_482;
  wire [7:0] coverage_36;
  wire  SaturatingCounter_73_clock;
  wire  SaturatingCounter_73_reset;
  wire  SaturatingCounter_73_io_enable;
  wire  SaturatingCounter_73_io_value;
  wire  _T_484;
  wire  SaturatingCounter_74_clock;
  wire  SaturatingCounter_74_reset;
  wire  SaturatingCounter_74_io_enable;
  wire  SaturatingCounter_74_io_value;
  wire  _T_485;
  wire [6:0] _T_489;
  wire [7:0] coverage_37;
  wire  SaturatingCounter_75_clock;
  wire  SaturatingCounter_75_reset;
  wire  SaturatingCounter_75_io_enable;
  wire  SaturatingCounter_75_io_value;
  wire  _T_491;
  wire  SaturatingCounter_76_clock;
  wire  SaturatingCounter_76_reset;
  wire  SaturatingCounter_76_io_enable;
  wire  SaturatingCounter_76_io_value;
  wire  _T_492;
  wire [6:0] _T_496;
  wire [7:0] coverage_38;
  wire  SaturatingCounter_77_clock;
  wire  SaturatingCounter_77_reset;
  wire  SaturatingCounter_77_io_enable;
  wire  SaturatingCounter_77_io_value;
  wire  _T_498;
  wire  SaturatingCounter_78_clock;
  wire  SaturatingCounter_78_reset;
  wire  SaturatingCounter_78_io_enable;
  wire  SaturatingCounter_78_io_value;
  wire  _T_499;
  wire [6:0] _T_503;
  wire [7:0] coverage_39;
  wire  SaturatingCounter_79_clock;
  wire  SaturatingCounter_79_reset;
  wire  SaturatingCounter_79_io_enable;
  wire  SaturatingCounter_79_io_value;
  wire  _T_505;
  wire  SaturatingCounter_80_clock;
  wire  SaturatingCounter_80_reset;
  wire  SaturatingCounter_80_io_enable;
  wire  SaturatingCounter_80_io_value;
  wire  _T_506;
  wire [6:0] _T_510;
  wire [7:0] coverage_40;
  wire  SaturatingCounter_81_clock;
  wire  SaturatingCounter_81_reset;
  wire  SaturatingCounter_81_io_enable;
  wire  SaturatingCounter_81_io_value;
  wire  _T_512;
  wire  SaturatingCounter_82_clock;
  wire  SaturatingCounter_82_reset;
  wire  SaturatingCounter_82_io_enable;
  wire  SaturatingCounter_82_io_value;
  wire  _T_513;
  wire [6:0] _T_517;
  wire [7:0] coverage_41;
  wire  SaturatingCounter_83_clock;
  wire  SaturatingCounter_83_reset;
  wire  SaturatingCounter_83_io_enable;
  wire  SaturatingCounter_83_io_value;
  wire  _T_519;
  wire  SaturatingCounter_84_clock;
  wire  SaturatingCounter_84_reset;
  wire  SaturatingCounter_84_io_enable;
  wire  SaturatingCounter_84_io_value;
  wire  _T_520;
  wire [6:0] _T_524;
  wire [7:0] coverage_42;
  wire  SaturatingCounter_85_clock;
  wire  SaturatingCounter_85_reset;
  wire  SaturatingCounter_85_io_enable;
  wire  SaturatingCounter_85_io_value;
  wire  _T_526;
  wire  SaturatingCounter_86_clock;
  wire  SaturatingCounter_86_reset;
  wire  SaturatingCounter_86_io_enable;
  wire  SaturatingCounter_86_io_value;
  wire  _T_527;
  wire [6:0] _T_531;
  wire [7:0] coverage_43;
  wire  SaturatingCounter_87_clock;
  wire  SaturatingCounter_87_reset;
  wire  SaturatingCounter_87_io_enable;
  wire  SaturatingCounter_87_io_value;
  wire  _T_533;
  wire  SaturatingCounter_88_clock;
  wire  SaturatingCounter_88_reset;
  wire  SaturatingCounter_88_io_enable;
  wire  SaturatingCounter_88_io_value;
  wire  _T_534;
  wire [6:0] _T_538;
  wire [7:0] coverage_44;
  wire  SaturatingCounter_89_clock;
  wire  SaturatingCounter_89_reset;
  wire  SaturatingCounter_89_io_enable;
  wire  SaturatingCounter_89_io_value;
  wire  _T_540;
  wire  SaturatingCounter_90_clock;
  wire  SaturatingCounter_90_reset;
  wire  SaturatingCounter_90_io_enable;
  wire  SaturatingCounter_90_io_value;
  wire  _T_541;
  wire [6:0] _T_545;
  wire [7:0] coverage_45;
  wire  SaturatingCounter_91_clock;
  wire  SaturatingCounter_91_reset;
  wire  SaturatingCounter_91_io_enable;
  wire  SaturatingCounter_91_io_value;
  wire  _T_547;
  wire  SaturatingCounter_92_clock;
  wire  SaturatingCounter_92_reset;
  wire  SaturatingCounter_92_io_enable;
  wire  SaturatingCounter_92_io_value;
  wire  _T_548;
  wire [6:0] _T_552;
  wire [7:0] coverage_46;
  wire  SaturatingCounter_93_clock;
  wire  SaturatingCounter_93_reset;
  wire  SaturatingCounter_93_io_enable;
  wire  SaturatingCounter_93_io_value;
  wire  _T_554;
  wire  SaturatingCounter_94_clock;
  wire  SaturatingCounter_94_reset;
  wire  SaturatingCounter_94_io_enable;
  wire  SaturatingCounter_94_io_value;
  wire  _T_555;
  wire [6:0] _T_559;
  wire [7:0] coverage_47;
  wire  SaturatingCounter_95_clock;
  wire  SaturatingCounter_95_reset;
  wire  SaturatingCounter_95_io_enable;
  wire  SaturatingCounter_95_io_value;
  wire  _T_561;
  wire  SaturatingCounter_96_clock;
  wire  SaturatingCounter_96_reset;
  wire  SaturatingCounter_96_io_enable;
  wire  SaturatingCounter_96_io_value;
  wire  _T_562;
  wire [6:0] _T_566;
  wire [7:0] coverage_48;
  wire  SaturatingCounter_97_clock;
  wire  SaturatingCounter_97_reset;
  wire  SaturatingCounter_97_io_enable;
  wire  SaturatingCounter_97_io_value;
  wire  _T_568;
  wire  SaturatingCounter_98_clock;
  wire  SaturatingCounter_98_reset;
  wire  SaturatingCounter_98_io_enable;
  wire  SaturatingCounter_98_io_value;
  wire  _T_569;
  wire [6:0] _T_573;
  wire [7:0] coverage_49;
  wire  SaturatingCounter_99_clock;
  wire  SaturatingCounter_99_reset;
  wire  SaturatingCounter_99_io_enable;
  wire  SaturatingCounter_99_io_value;
  wire  _T_575;
  wire  SaturatingCounter_100_clock;
  wire  SaturatingCounter_100_reset;
  wire  SaturatingCounter_100_io_enable;
  wire  SaturatingCounter_100_io_value;
  wire  _T_576;
  wire [6:0] _T_580;
  wire [7:0] coverage_50;
  wire  SaturatingCounter_101_clock;
  wire  SaturatingCounter_101_reset;
  wire  SaturatingCounter_101_io_enable;
  wire  SaturatingCounter_101_io_value;
  wire  _T_582;
  wire  SaturatingCounter_102_clock;
  wire  SaturatingCounter_102_reset;
  wire  SaturatingCounter_102_io_enable;
  wire  SaturatingCounter_102_io_value;
  wire  _T_583;
  wire [6:0] _T_587;
  wire [7:0] coverage_51;
  wire  SaturatingCounter_103_clock;
  wire  SaturatingCounter_103_reset;
  wire  SaturatingCounter_103_io_enable;
  wire  SaturatingCounter_103_io_value;
  wire  _T_589;
  wire  SaturatingCounter_104_clock;
  wire  SaturatingCounter_104_reset;
  wire  SaturatingCounter_104_io_enable;
  wire  SaturatingCounter_104_io_value;
  wire  _T_590;
  wire [6:0] _T_594;
  wire [7:0] coverage_52;
  wire  SaturatingCounter_105_clock;
  wire  SaturatingCounter_105_reset;
  wire  SaturatingCounter_105_io_enable;
  wire  SaturatingCounter_105_io_value;
  wire  _T_596;
  wire  SaturatingCounter_106_clock;
  wire  SaturatingCounter_106_reset;
  wire  SaturatingCounter_106_io_enable;
  wire  SaturatingCounter_106_io_value;
  wire  _T_597;
  wire [6:0] _T_601;
  wire [7:0] coverage_53;
  wire  SaturatingCounter_107_clock;
  wire  SaturatingCounter_107_reset;
  wire  SaturatingCounter_107_io_enable;
  wire  SaturatingCounter_107_io_value;
  wire  _T_603;
  wire  SaturatingCounter_108_clock;
  wire  SaturatingCounter_108_reset;
  wire  SaturatingCounter_108_io_enable;
  wire  SaturatingCounter_108_io_value;
  wire  _T_604;
  wire [6:0] _T_608;
  wire [7:0] coverage_54;
  wire  SaturatingCounter_109_clock;
  wire  SaturatingCounter_109_reset;
  wire  SaturatingCounter_109_io_enable;
  wire  SaturatingCounter_109_io_value;
  wire  _T_610;
  wire  SaturatingCounter_110_clock;
  wire  SaturatingCounter_110_reset;
  wire  SaturatingCounter_110_io_enable;
  wire  SaturatingCounter_110_io_value;
  wire  _T_611;
  wire [6:0] _T_615;
  wire [7:0] coverage_55;
  wire  SaturatingCounter_111_clock;
  wire  SaturatingCounter_111_reset;
  wire  SaturatingCounter_111_io_enable;
  wire  SaturatingCounter_111_io_value;
  wire  _T_617;
  wire  SaturatingCounter_112_clock;
  wire  SaturatingCounter_112_reset;
  wire  SaturatingCounter_112_io_enable;
  wire  SaturatingCounter_112_io_value;
  wire  _T_618;
  wire [6:0] _T_622;
  wire [7:0] coverage_56;
  wire  SaturatingCounter_113_clock;
  wire  SaturatingCounter_113_reset;
  wire  SaturatingCounter_113_io_enable;
  wire  SaturatingCounter_113_io_value;
  wire  _T_624;
  wire  SaturatingCounter_114_clock;
  wire  SaturatingCounter_114_reset;
  wire  SaturatingCounter_114_io_enable;
  wire  SaturatingCounter_114_io_value;
  wire  _T_625;
  wire [6:0] _T_629;
  wire [7:0] coverage_57;
  wire  SaturatingCounter_115_clock;
  wire  SaturatingCounter_115_reset;
  wire  SaturatingCounter_115_io_enable;
  wire  SaturatingCounter_115_io_value;
  wire  _T_631;
  wire  SaturatingCounter_116_clock;
  wire  SaturatingCounter_116_reset;
  wire  SaturatingCounter_116_io_enable;
  wire  SaturatingCounter_116_io_value;
  wire  _T_632;
  wire [6:0] _T_636;
  wire [7:0] coverage_58;
  wire  SaturatingCounter_117_clock;
  wire  SaturatingCounter_117_reset;
  wire  SaturatingCounter_117_io_enable;
  wire  SaturatingCounter_117_io_value;
  wire  _T_638;
  wire  SaturatingCounter_118_clock;
  wire  SaturatingCounter_118_reset;
  wire  SaturatingCounter_118_io_enable;
  wire  SaturatingCounter_118_io_value;
  wire  _T_639;
  wire [6:0] _T_643;
  wire [7:0] coverage_59;
  wire  SaturatingCounter_119_clock;
  wire  SaturatingCounter_119_reset;
  wire  SaturatingCounter_119_io_enable;
  wire  SaturatingCounter_119_io_value;
  wire  _T_645;
  wire  SaturatingCounter_120_clock;
  wire  SaturatingCounter_120_reset;
  wire  SaturatingCounter_120_io_enable;
  wire  SaturatingCounter_120_io_value;
  wire  _T_646;
  wire [6:0] _T_650;
  wire [7:0] coverage_60;
  wire  SaturatingCounter_121_clock;
  wire  SaturatingCounter_121_reset;
  wire  SaturatingCounter_121_io_enable;
  wire  SaturatingCounter_121_io_value;
  wire  _T_652;
  wire  SaturatingCounter_122_clock;
  wire  SaturatingCounter_122_reset;
  wire  SaturatingCounter_122_io_enable;
  wire  SaturatingCounter_122_io_value;
  wire  _T_653;
  wire [6:0] _T_657;
  wire [7:0] coverage_61;
  wire  SaturatingCounter_123_clock;
  wire  SaturatingCounter_123_reset;
  wire  SaturatingCounter_123_io_enable;
  wire  SaturatingCounter_123_io_value;
  wire  _T_659;
  wire  SaturatingCounter_124_clock;
  wire  SaturatingCounter_124_reset;
  wire  SaturatingCounter_124_io_enable;
  wire  SaturatingCounter_124_io_value;
  wire  _T_660;
  wire [6:0] _T_664;
  wire [7:0] coverage_62;
  wire  SaturatingCounter_125_clock;
  wire  SaturatingCounter_125_reset;
  wire  SaturatingCounter_125_io_enable;
  wire  SaturatingCounter_125_io_value;
  wire  _T_666;
  wire  SaturatingCounter_126_clock;
  wire  SaturatingCounter_126_reset;
  wire  SaturatingCounter_126_io_enable;
  wire  SaturatingCounter_126_io_value;
  wire  _T_667;
  wire [6:0] _T_671;
  wire [7:0] coverage_63;
  wire  SaturatingCounter_127_clock;
  wire  SaturatingCounter_127_reset;
  wire  SaturatingCounter_127_io_enable;
  wire  SaturatingCounter_127_io_value;
  wire  _T_673;
  wire  SaturatingCounter_128_clock;
  wire  SaturatingCounter_128_reset;
  wire  SaturatingCounter_128_io_enable;
  wire  SaturatingCounter_128_io_value;
  wire  _T_674;
  wire [6:0] _T_678;
  wire [7:0] coverage_64;
  wire  SaturatingCounter_129_clock;
  wire  SaturatingCounter_129_reset;
  wire  SaturatingCounter_129_io_enable;
  wire  SaturatingCounter_129_io_value;
  wire  _T_680;
  wire  SaturatingCounter_130_clock;
  wire  SaturatingCounter_130_reset;
  wire  SaturatingCounter_130_io_enable;
  wire  SaturatingCounter_130_io_value;
  wire  _T_681;
  wire [6:0] _T_685;
  wire [7:0] coverage_65;
  wire  SaturatingCounter_131_clock;
  wire  SaturatingCounter_131_reset;
  wire  SaturatingCounter_131_io_enable;
  wire  SaturatingCounter_131_io_value;
  wire  _T_687;
  wire  SaturatingCounter_132_clock;
  wire  SaturatingCounter_132_reset;
  wire  SaturatingCounter_132_io_enable;
  wire  SaturatingCounter_132_io_value;
  wire  _T_688;
  wire [6:0] _T_692;
  wire [7:0] coverage_66;
  wire  SaturatingCounter_133_clock;
  wire  SaturatingCounter_133_reset;
  wire  SaturatingCounter_133_io_enable;
  wire  SaturatingCounter_133_io_value;
  wire  _T_694;
  wire  SaturatingCounter_134_clock;
  wire  SaturatingCounter_134_reset;
  wire  SaturatingCounter_134_io_enable;
  wire  SaturatingCounter_134_io_value;
  wire  _T_695;
  wire [6:0] _T_699;
  wire [7:0] coverage_67;
  wire  SaturatingCounter_135_clock;
  wire  SaturatingCounter_135_reset;
  wire  SaturatingCounter_135_io_enable;
  wire  SaturatingCounter_135_io_value;
  wire  _T_701;
  wire  SaturatingCounter_136_clock;
  wire  SaturatingCounter_136_reset;
  wire  SaturatingCounter_136_io_enable;
  wire  SaturatingCounter_136_io_value;
  wire  _T_702;
  wire [6:0] _T_706;
  wire [7:0] coverage_68;
  wire  SaturatingCounter_137_clock;
  wire  SaturatingCounter_137_reset;
  wire  SaturatingCounter_137_io_enable;
  wire  SaturatingCounter_137_io_value;
  wire  _T_708;
  wire  SaturatingCounter_138_clock;
  wire  SaturatingCounter_138_reset;
  wire  SaturatingCounter_138_io_enable;
  wire  SaturatingCounter_138_io_value;
  wire  _T_709;
  wire [6:0] _T_713;
  wire [7:0] coverage_69;
  wire  SaturatingCounter_139_clock;
  wire  SaturatingCounter_139_reset;
  wire  SaturatingCounter_139_io_enable;
  wire  SaturatingCounter_139_io_value;
  wire  _T_715;
  wire  SaturatingCounter_140_clock;
  wire  SaturatingCounter_140_reset;
  wire  SaturatingCounter_140_io_enable;
  wire  SaturatingCounter_140_io_value;
  wire  _T_716;
  wire [6:0] _T_720;
  wire [7:0] coverage_70;
  wire  SaturatingCounter_141_clock;
  wire  SaturatingCounter_141_reset;
  wire  SaturatingCounter_141_io_enable;
  wire  SaturatingCounter_141_io_value;
  wire  _T_722;
  wire  SaturatingCounter_142_clock;
  wire  SaturatingCounter_142_reset;
  wire  SaturatingCounter_142_io_enable;
  wire  SaturatingCounter_142_io_value;
  wire  _T_723;
  wire [6:0] _T_727;
  wire [7:0] coverage_71;
  wire  SaturatingCounter_143_clock;
  wire  SaturatingCounter_143_reset;
  wire  SaturatingCounter_143_io_enable;
  wire  SaturatingCounter_143_io_value;
  wire  _T_729;
  wire  SaturatingCounter_144_clock;
  wire  SaturatingCounter_144_reset;
  wire  SaturatingCounter_144_io_enable;
  wire  SaturatingCounter_144_io_value;
  wire  _T_730;
  wire [6:0] _T_734;
  wire [7:0] coverage_72;
  wire  SaturatingCounter_145_clock;
  wire  SaturatingCounter_145_reset;
  wire  SaturatingCounter_145_io_enable;
  wire  SaturatingCounter_145_io_value;
  wire  _T_736;
  wire  SaturatingCounter_146_clock;
  wire  SaturatingCounter_146_reset;
  wire  SaturatingCounter_146_io_enable;
  wire  SaturatingCounter_146_io_value;
  wire  _T_737;
  wire [6:0] _T_741;
  wire [7:0] coverage_73;
  wire  SaturatingCounter_147_clock;
  wire  SaturatingCounter_147_reset;
  wire  SaturatingCounter_147_io_enable;
  wire  SaturatingCounter_147_io_value;
  wire  _T_743;
  wire  SaturatingCounter_148_clock;
  wire  SaturatingCounter_148_reset;
  wire  SaturatingCounter_148_io_enable;
  wire  SaturatingCounter_148_io_value;
  wire  _T_744;
  wire [6:0] _T_748;
  wire [7:0] coverage_74;
  wire  SaturatingCounter_149_clock;
  wire  SaturatingCounter_149_reset;
  wire  SaturatingCounter_149_io_enable;
  wire  SaturatingCounter_149_io_value;
  wire  _T_750;
  wire  SaturatingCounter_150_clock;
  wire  SaturatingCounter_150_reset;
  wire  SaturatingCounter_150_io_enable;
  wire  SaturatingCounter_150_io_value;
  wire  _T_751;
  wire [6:0] _T_755;
  wire [7:0] coverage_75;
  wire  SaturatingCounter_151_clock;
  wire  SaturatingCounter_151_reset;
  wire  SaturatingCounter_151_io_enable;
  wire  SaturatingCounter_151_io_value;
  wire  _T_757;
  wire  SaturatingCounter_152_clock;
  wire  SaturatingCounter_152_reset;
  wire  SaturatingCounter_152_io_enable;
  wire  SaturatingCounter_152_io_value;
  wire  _T_758;
  wire [6:0] _T_762;
  wire [7:0] coverage_76;
  wire  SaturatingCounter_153_clock;
  wire  SaturatingCounter_153_reset;
  wire  SaturatingCounter_153_io_enable;
  wire  SaturatingCounter_153_io_value;
  wire  _T_764;
  wire  SaturatingCounter_154_clock;
  wire  SaturatingCounter_154_reset;
  wire  SaturatingCounter_154_io_enable;
  wire  SaturatingCounter_154_io_value;
  wire  _T_765;
  wire [6:0] _T_769;
  wire [7:0] coverage_77;
  wire  SaturatingCounter_155_clock;
  wire  SaturatingCounter_155_reset;
  wire  SaturatingCounter_155_io_enable;
  wire  SaturatingCounter_155_io_value;
  wire  _T_771;
  wire  SaturatingCounter_156_clock;
  wire  SaturatingCounter_156_reset;
  wire  SaturatingCounter_156_io_enable;
  wire  SaturatingCounter_156_io_value;
  wire  _T_772;
  wire [6:0] _T_776;
  wire [7:0] coverage_78;
  wire  SaturatingCounter_157_clock;
  wire  SaturatingCounter_157_reset;
  wire  SaturatingCounter_157_io_enable;
  wire  SaturatingCounter_157_io_value;
  wire  _T_778;
  wire  SaturatingCounter_158_clock;
  wire  SaturatingCounter_158_reset;
  wire  SaturatingCounter_158_io_enable;
  wire  SaturatingCounter_158_io_value;
  wire  _T_779;
  wire [6:0] _T_783;
  wire [7:0] coverage_79;
  wire  SaturatingCounter_159_clock;
  wire  SaturatingCounter_159_reset;
  wire  SaturatingCounter_159_io_enable;
  wire  SaturatingCounter_159_io_value;
  wire  _T_785;
  wire  SaturatingCounter_160_clock;
  wire  SaturatingCounter_160_reset;
  wire  SaturatingCounter_160_io_enable;
  wire  SaturatingCounter_160_io_value;
  wire  _T_786;
  wire [6:0] _T_790;
  wire [7:0] coverage_80;
  wire  SaturatingCounter_161_clock;
  wire  SaturatingCounter_161_reset;
  wire  SaturatingCounter_161_io_enable;
  wire  SaturatingCounter_161_io_value;
  wire  _T_792;
  wire  SaturatingCounter_162_clock;
  wire  SaturatingCounter_162_reset;
  wire  SaturatingCounter_162_io_enable;
  wire  SaturatingCounter_162_io_value;
  wire  _T_793;
  wire [6:0] _T_797;
  wire [7:0] coverage_81;
  wire  SaturatingCounter_163_clock;
  wire  SaturatingCounter_163_reset;
  wire  SaturatingCounter_163_io_enable;
  wire  SaturatingCounter_163_io_value;
  wire  _T_799;
  wire  SaturatingCounter_164_clock;
  wire  SaturatingCounter_164_reset;
  wire  SaturatingCounter_164_io_enable;
  wire  SaturatingCounter_164_io_value;
  wire  _T_800;
  wire [6:0] _T_804;
  wire [7:0] coverage_82;
  wire  SaturatingCounter_165_clock;
  wire  SaturatingCounter_165_reset;
  wire  SaturatingCounter_165_io_enable;
  wire  SaturatingCounter_165_io_value;
  wire  _T_806;
  wire  SaturatingCounter_166_clock;
  wire  SaturatingCounter_166_reset;
  wire  SaturatingCounter_166_io_enable;
  wire  SaturatingCounter_166_io_value;
  wire  _T_807;
  wire [6:0] _T_811;
  wire [7:0] coverage_83;
  wire  SaturatingCounter_167_clock;
  wire  SaturatingCounter_167_reset;
  wire  SaturatingCounter_167_io_enable;
  wire  SaturatingCounter_167_io_value;
  wire  _T_813;
  wire  SaturatingCounter_168_clock;
  wire  SaturatingCounter_168_reset;
  wire  SaturatingCounter_168_io_enable;
  wire  SaturatingCounter_168_io_value;
  wire  _T_814;
  wire [6:0] _T_818;
  wire [7:0] coverage_84;
  wire  SaturatingCounter_169_clock;
  wire  SaturatingCounter_169_reset;
  wire  SaturatingCounter_169_io_enable;
  wire  SaturatingCounter_169_io_value;
  wire  _T_820;
  wire  SaturatingCounter_170_clock;
  wire  SaturatingCounter_170_reset;
  wire  SaturatingCounter_170_io_enable;
  wire  SaturatingCounter_170_io_value;
  wire  _T_821;
  wire [6:0] _T_825;
  wire [7:0] coverage_85;
  wire  SaturatingCounter_171_clock;
  wire  SaturatingCounter_171_reset;
  wire  SaturatingCounter_171_io_enable;
  wire  SaturatingCounter_171_io_value;
  wire  _T_827;
  wire  SaturatingCounter_172_clock;
  wire  SaturatingCounter_172_reset;
  wire  SaturatingCounter_172_io_enable;
  wire  SaturatingCounter_172_io_value;
  wire  _T_828;
  wire [6:0] _T_832;
  wire [7:0] coverage_86;
  wire  SaturatingCounter_173_clock;
  wire  SaturatingCounter_173_reset;
  wire  SaturatingCounter_173_io_enable;
  wire  SaturatingCounter_173_io_value;
  wire  _T_834;
  wire  SaturatingCounter_174_clock;
  wire  SaturatingCounter_174_reset;
  wire  SaturatingCounter_174_io_enable;
  wire  SaturatingCounter_174_io_value;
  wire  _T_835;
  wire [6:0] _T_839;
  wire [7:0] coverage_87;
  wire  SaturatingCounter_175_clock;
  wire  SaturatingCounter_175_reset;
  wire  SaturatingCounter_175_io_enable;
  wire  SaturatingCounter_175_io_value;
  wire  _T_841;
  wire  SaturatingCounter_176_clock;
  wire  SaturatingCounter_176_reset;
  wire  SaturatingCounter_176_io_enable;
  wire  SaturatingCounter_176_io_value;
  wire  _T_842;
  wire [6:0] _T_846;
  wire [7:0] coverage_88;
  wire  SaturatingCounter_177_clock;
  wire  SaturatingCounter_177_reset;
  wire  SaturatingCounter_177_io_enable;
  wire  SaturatingCounter_177_io_value;
  wire  _T_848;
  wire  SaturatingCounter_178_clock;
  wire  SaturatingCounter_178_reset;
  wire  SaturatingCounter_178_io_enable;
  wire  SaturatingCounter_178_io_value;
  wire  _T_849;
  wire [6:0] _T_853;
  wire [7:0] coverage_89;
  wire  SaturatingCounter_179_clock;
  wire  SaturatingCounter_179_reset;
  wire  SaturatingCounter_179_io_enable;
  wire  SaturatingCounter_179_io_value;
  wire  _T_855;
  wire  SaturatingCounter_180_clock;
  wire  SaturatingCounter_180_reset;
  wire  SaturatingCounter_180_io_enable;
  wire  SaturatingCounter_180_io_value;
  wire  _T_856;
  wire [6:0] _T_860;
  wire [7:0] coverage_90;
  wire  SaturatingCounter_181_clock;
  wire  SaturatingCounter_181_reset;
  wire  SaturatingCounter_181_io_enable;
  wire  SaturatingCounter_181_io_value;
  wire  _T_862;
  wire  SaturatingCounter_182_clock;
  wire  SaturatingCounter_182_reset;
  wire  SaturatingCounter_182_io_enable;
  wire  SaturatingCounter_182_io_value;
  wire  _T_863;
  wire [6:0] _T_867;
  wire [7:0] coverage_91;
  wire  SaturatingCounter_183_clock;
  wire  SaturatingCounter_183_reset;
  wire  SaturatingCounter_183_io_enable;
  wire  SaturatingCounter_183_io_value;
  wire  _T_869;
  wire  SaturatingCounter_184_clock;
  wire  SaturatingCounter_184_reset;
  wire  SaturatingCounter_184_io_enable;
  wire  SaturatingCounter_184_io_value;
  wire  _T_870;
  wire [6:0] _T_874;
  wire [7:0] coverage_92;
  wire  SaturatingCounter_185_clock;
  wire  SaturatingCounter_185_reset;
  wire  SaturatingCounter_185_io_enable;
  wire  SaturatingCounter_185_io_value;
  wire  _T_876;
  wire  SaturatingCounter_186_clock;
  wire  SaturatingCounter_186_reset;
  wire  SaturatingCounter_186_io_enable;
  wire  SaturatingCounter_186_io_value;
  wire  _T_877;
  wire [6:0] _T_881;
  wire [7:0] coverage_93;
  wire  SaturatingCounter_187_clock;
  wire  SaturatingCounter_187_reset;
  wire  SaturatingCounter_187_io_enable;
  wire  SaturatingCounter_187_io_value;
  wire  _T_883;
  wire  SaturatingCounter_188_clock;
  wire  SaturatingCounter_188_reset;
  wire  SaturatingCounter_188_io_enable;
  wire  SaturatingCounter_188_io_value;
  wire  _T_884;
  wire [6:0] _T_888;
  wire [7:0] coverage_94;
  wire  SaturatingCounter_189_clock;
  wire  SaturatingCounter_189_reset;
  wire  SaturatingCounter_189_io_enable;
  wire  SaturatingCounter_189_io_value;
  wire  _T_890;
  wire  SaturatingCounter_190_clock;
  wire  SaturatingCounter_190_reset;
  wire  SaturatingCounter_190_io_enable;
  wire  SaturatingCounter_190_io_value;
  wire  _T_891;
  wire [6:0] _T_895;
  wire [7:0] coverage_95;
  wire  SaturatingCounter_191_clock;
  wire  SaturatingCounter_191_reset;
  wire  SaturatingCounter_191_io_enable;
  wire  SaturatingCounter_191_io_value;
  wire  _T_897;
  wire  SaturatingCounter_192_clock;
  wire  SaturatingCounter_192_reset;
  wire  SaturatingCounter_192_io_enable;
  wire  SaturatingCounter_192_io_value;
  wire  _T_898;
  wire [6:0] _T_902;
  wire [7:0] coverage_96;
  wire  SaturatingCounter_193_clock;
  wire  SaturatingCounter_193_reset;
  wire  SaturatingCounter_193_io_enable;
  wire  SaturatingCounter_193_io_value;
  wire  _T_904;
  wire  SaturatingCounter_194_clock;
  wire  SaturatingCounter_194_reset;
  wire  SaturatingCounter_194_io_enable;
  wire  SaturatingCounter_194_io_value;
  wire  _T_905;
  wire [6:0] _T_909;
  wire [7:0] coverage_97;
  wire  SaturatingCounter_195_clock;
  wire  SaturatingCounter_195_reset;
  wire  SaturatingCounter_195_io_enable;
  wire  SaturatingCounter_195_io_value;
  wire  _T_911;
  wire  SaturatingCounter_196_clock;
  wire  SaturatingCounter_196_reset;
  wire  SaturatingCounter_196_io_enable;
  wire  SaturatingCounter_196_io_value;
  wire  _T_912;
  wire [6:0] _T_916;
  wire [7:0] coverage_98;
  wire  SaturatingCounter_197_clock;
  wire  SaturatingCounter_197_reset;
  wire  SaturatingCounter_197_io_enable;
  wire  SaturatingCounter_197_io_value;
  wire  _T_918;
  wire  SaturatingCounter_198_clock;
  wire  SaturatingCounter_198_reset;
  wire  SaturatingCounter_198_io_enable;
  wire  SaturatingCounter_198_io_value;
  wire  _T_919;
  wire [6:0] _T_923;
  wire [7:0] coverage_99;
  wire  SaturatingCounter_199_clock;
  wire  SaturatingCounter_199_reset;
  wire  SaturatingCounter_199_io_enable;
  wire  SaturatingCounter_199_io_value;
  wire  _T_925;
  wire  SaturatingCounter_200_clock;
  wire  SaturatingCounter_200_reset;
  wire  SaturatingCounter_200_io_enable;
  wire  SaturatingCounter_200_io_value;
  wire  _T_926;
  wire [6:0] _T_930;
  wire [7:0] coverage_100;
  wire  SaturatingCounter_201_clock;
  wire  SaturatingCounter_201_reset;
  wire  SaturatingCounter_201_io_enable;
  wire  SaturatingCounter_201_io_value;
  wire  _T_932;
  wire  SaturatingCounter_202_clock;
  wire  SaturatingCounter_202_reset;
  wire  SaturatingCounter_202_io_enable;
  wire  SaturatingCounter_202_io_value;
  wire  _T_933;
  wire [6:0] _T_937;
  wire [7:0] coverage_101;
  wire  SaturatingCounter_203_clock;
  wire  SaturatingCounter_203_reset;
  wire  SaturatingCounter_203_io_enable;
  wire  SaturatingCounter_203_io_value;
  wire  _T_939;
  wire  SaturatingCounter_204_clock;
  wire  SaturatingCounter_204_reset;
  wire  SaturatingCounter_204_io_enable;
  wire  SaturatingCounter_204_io_value;
  wire  _T_940;
  wire [6:0] _T_944;
  wire [7:0] coverage_102;
  wire  SaturatingCounter_205_clock;
  wire  SaturatingCounter_205_reset;
  wire  SaturatingCounter_205_io_enable;
  wire  SaturatingCounter_205_io_value;
  wire  _T_946;
  wire  SaturatingCounter_206_clock;
  wire  SaturatingCounter_206_reset;
  wire  SaturatingCounter_206_io_enable;
  wire  SaturatingCounter_206_io_value;
  wire  _T_947;
  wire [6:0] _T_951;
  wire [7:0] coverage_103;
  wire  SaturatingCounter_207_clock;
  wire  SaturatingCounter_207_reset;
  wire  SaturatingCounter_207_io_enable;
  wire  SaturatingCounter_207_io_value;
  wire  _T_953;
  wire  SaturatingCounter_208_clock;
  wire  SaturatingCounter_208_reset;
  wire  SaturatingCounter_208_io_enable;
  wire  SaturatingCounter_208_io_value;
  wire  _T_954;
  wire [6:0] _T_958;
  wire [7:0] coverage_104;
  wire  SaturatingCounter_209_clock;
  wire  SaturatingCounter_209_reset;
  wire  SaturatingCounter_209_io_enable;
  wire  SaturatingCounter_209_io_value;
  wire  _T_960;
  wire  SaturatingCounter_210_clock;
  wire  SaturatingCounter_210_reset;
  wire  SaturatingCounter_210_io_enable;
  wire  SaturatingCounter_210_io_value;
  wire  _T_961;
  wire [6:0] _T_965;
  wire [7:0] coverage_105;
  wire  SaturatingCounter_211_clock;
  wire  SaturatingCounter_211_reset;
  wire  SaturatingCounter_211_io_enable;
  wire  SaturatingCounter_211_io_value;
  wire  _T_967;
  wire  SaturatingCounter_212_clock;
  wire  SaturatingCounter_212_reset;
  wire  SaturatingCounter_212_io_enable;
  wire  SaturatingCounter_212_io_value;
  wire  _T_968;
  wire [6:0] _T_972;
  wire [7:0] coverage_106;
  wire  SaturatingCounter_213_clock;
  wire  SaturatingCounter_213_reset;
  wire  SaturatingCounter_213_io_enable;
  wire  SaturatingCounter_213_io_value;
  wire  _T_974;
  wire  SaturatingCounter_214_clock;
  wire  SaturatingCounter_214_reset;
  wire  SaturatingCounter_214_io_enable;
  wire  SaturatingCounter_214_io_value;
  wire  _T_975;
  wire [6:0] _T_979;
  wire [7:0] coverage_107;
  wire  SaturatingCounter_215_clock;
  wire  SaturatingCounter_215_reset;
  wire  SaturatingCounter_215_io_enable;
  wire  SaturatingCounter_215_io_value;
  wire  _T_981;
  wire  SaturatingCounter_216_clock;
  wire  SaturatingCounter_216_reset;
  wire  SaturatingCounter_216_io_enable;
  wire  SaturatingCounter_216_io_value;
  wire  _T_982;
  wire [6:0] _T_986;
  wire [7:0] coverage_108;
  wire  SaturatingCounter_217_clock;
  wire  SaturatingCounter_217_reset;
  wire  SaturatingCounter_217_io_enable;
  wire  SaturatingCounter_217_io_value;
  wire  _T_988;
  wire  SaturatingCounter_218_clock;
  wire  SaturatingCounter_218_reset;
  wire  SaturatingCounter_218_io_enable;
  wire  SaturatingCounter_218_io_value;
  wire  _T_989;
  wire [6:0] _T_993;
  wire [7:0] coverage_109;
  wire  SaturatingCounter_219_clock;
  wire  SaturatingCounter_219_reset;
  wire  SaturatingCounter_219_io_enable;
  wire  SaturatingCounter_219_io_value;
  wire  _T_995;
  wire  SaturatingCounter_220_clock;
  wire  SaturatingCounter_220_reset;
  wire  SaturatingCounter_220_io_enable;
  wire  SaturatingCounter_220_io_value;
  wire  _T_996;
  wire [6:0] _T_1000;
  wire [7:0] coverage_110;
  wire  SaturatingCounter_221_clock;
  wire  SaturatingCounter_221_reset;
  wire  SaturatingCounter_221_io_enable;
  wire  SaturatingCounter_221_io_value;
  wire  _T_1002;
  wire  SaturatingCounter_222_clock;
  wire  SaturatingCounter_222_reset;
  wire  SaturatingCounter_222_io_enable;
  wire  SaturatingCounter_222_io_value;
  wire  _T_1003;
  wire [6:0] _T_1007;
  wire [7:0] coverage_111;
  wire  SaturatingCounter_223_clock;
  wire  SaturatingCounter_223_reset;
  wire  SaturatingCounter_223_io_enable;
  wire  SaturatingCounter_223_io_value;
  wire  _T_1009;
  wire  SaturatingCounter_224_clock;
  wire  SaturatingCounter_224_reset;
  wire  SaturatingCounter_224_io_enable;
  wire  SaturatingCounter_224_io_value;
  wire  _T_1010;
  wire [6:0] _T_1014;
  wire [7:0] coverage_112;
  wire  SaturatingCounter_225_clock;
  wire  SaturatingCounter_225_reset;
  wire  SaturatingCounter_225_io_enable;
  wire  SaturatingCounter_225_io_value;
  wire  _T_1016;
  wire  SaturatingCounter_226_clock;
  wire  SaturatingCounter_226_reset;
  wire  SaturatingCounter_226_io_enable;
  wire  SaturatingCounter_226_io_value;
  wire  _T_1017;
  wire [6:0] _T_1021;
  wire [7:0] coverage_113;
  wire  SaturatingCounter_227_clock;
  wire  SaturatingCounter_227_reset;
  wire  SaturatingCounter_227_io_enable;
  wire  SaturatingCounter_227_io_value;
  wire  _T_1023;
  wire  SaturatingCounter_228_clock;
  wire  SaturatingCounter_228_reset;
  wire  SaturatingCounter_228_io_enable;
  wire  SaturatingCounter_228_io_value;
  wire  _T_1024;
  wire [6:0] _T_1028;
  wire [7:0] coverage_114;
  wire  SaturatingCounter_229_clock;
  wire  SaturatingCounter_229_reset;
  wire  SaturatingCounter_229_io_enable;
  wire  SaturatingCounter_229_io_value;
  wire  _T_1030;
  wire  SaturatingCounter_230_clock;
  wire  SaturatingCounter_230_reset;
  wire  SaturatingCounter_230_io_enable;
  wire  SaturatingCounter_230_io_value;
  wire  _T_1031;
  wire [6:0] _T_1035;
  wire [7:0] coverage_115;
  wire  SaturatingCounter_231_clock;
  wire  SaturatingCounter_231_reset;
  wire  SaturatingCounter_231_io_enable;
  wire  SaturatingCounter_231_io_value;
  wire  _T_1037;
  wire  SaturatingCounter_232_clock;
  wire  SaturatingCounter_232_reset;
  wire  SaturatingCounter_232_io_enable;
  wire  SaturatingCounter_232_io_value;
  wire  _T_1038;
  wire [6:0] _T_1042;
  wire [7:0] coverage_116;
  wire  SaturatingCounter_233_clock;
  wire  SaturatingCounter_233_reset;
  wire  SaturatingCounter_233_io_enable;
  wire  SaturatingCounter_233_io_value;
  wire  _T_1044;
  wire  SaturatingCounter_234_clock;
  wire  SaturatingCounter_234_reset;
  wire  SaturatingCounter_234_io_enable;
  wire  SaturatingCounter_234_io_value;
  wire  _T_1045;
  wire [6:0] _T_1049;
  wire [7:0] coverage_117;
  wire  SaturatingCounter_235_clock;
  wire  SaturatingCounter_235_reset;
  wire  SaturatingCounter_235_io_enable;
  wire  SaturatingCounter_235_io_value;
  wire  _T_1051;
  wire  SaturatingCounter_236_clock;
  wire  SaturatingCounter_236_reset;
  wire  SaturatingCounter_236_io_enable;
  wire  SaturatingCounter_236_io_value;
  wire  _T_1052;
  wire [6:0] _T_1056;
  wire [7:0] coverage_118;
  wire  SaturatingCounter_237_clock;
  wire  SaturatingCounter_237_reset;
  wire  SaturatingCounter_237_io_enable;
  wire  SaturatingCounter_237_io_value;
  wire  _T_1058;
  wire  SaturatingCounter_238_clock;
  wire  SaturatingCounter_238_reset;
  wire  SaturatingCounter_238_io_enable;
  wire  SaturatingCounter_238_io_value;
  wire  _T_1059;
  wire [6:0] _T_1063;
  wire [7:0] coverage_119;
  wire  SaturatingCounter_239_clock;
  wire  SaturatingCounter_239_reset;
  wire  SaturatingCounter_239_io_enable;
  wire  SaturatingCounter_239_io_value;
  wire  _T_1065;
  wire  SaturatingCounter_240_clock;
  wire  SaturatingCounter_240_reset;
  wire  SaturatingCounter_240_io_enable;
  wire  SaturatingCounter_240_io_value;
  wire  _T_1066;
  wire [6:0] _T_1070;
  wire [7:0] coverage_120;
  wire  SaturatingCounter_241_clock;
  wire  SaturatingCounter_241_reset;
  wire  SaturatingCounter_241_io_enable;
  wire  SaturatingCounter_241_io_value;
  wire  _T_1072;
  wire  SaturatingCounter_242_clock;
  wire  SaturatingCounter_242_reset;
  wire  SaturatingCounter_242_io_enable;
  wire  SaturatingCounter_242_io_value;
  wire  _T_1073;
  wire [6:0] _T_1077;
  wire [7:0] coverage_121;
  wire  SaturatingCounter_243_clock;
  wire  SaturatingCounter_243_reset;
  wire  SaturatingCounter_243_io_enable;
  wire  SaturatingCounter_243_io_value;
  wire  _T_1079;
  wire  SaturatingCounter_244_clock;
  wire  SaturatingCounter_244_reset;
  wire  SaturatingCounter_244_io_enable;
  wire  SaturatingCounter_244_io_value;
  wire  _T_1080;
  wire [6:0] _T_1084;
  wire [7:0] coverage_122;
  wire  SaturatingCounter_245_clock;
  wire  SaturatingCounter_245_reset;
  wire  SaturatingCounter_245_io_enable;
  wire  SaturatingCounter_245_io_value;
  wire  _T_1086;
  wire  SaturatingCounter_246_clock;
  wire  SaturatingCounter_246_reset;
  wire  SaturatingCounter_246_io_enable;
  wire  SaturatingCounter_246_io_value;
  wire  _T_1087;
  wire [6:0] _T_1091;
  wire [7:0] coverage_123;
  wire  SaturatingCounter_247_clock;
  wire  SaturatingCounter_247_reset;
  wire  SaturatingCounter_247_io_enable;
  wire  SaturatingCounter_247_io_value;
  wire  _T_1093;
  wire  SaturatingCounter_248_clock;
  wire  SaturatingCounter_248_reset;
  wire  SaturatingCounter_248_io_enable;
  wire  SaturatingCounter_248_io_value;
  wire  _T_1094;
  wire [6:0] _T_1098;
  wire [7:0] coverage_124;
  wire  SaturatingCounter_249_clock;
  wire  SaturatingCounter_249_reset;
  wire  SaturatingCounter_249_io_enable;
  wire  SaturatingCounter_249_io_value;
  wire  _T_1100;
  wire  SaturatingCounter_250_clock;
  wire  SaturatingCounter_250_reset;
  wire  SaturatingCounter_250_io_enable;
  wire  SaturatingCounter_250_io_value;
  wire  _T_1101;
  wire [6:0] _T_1105;
  wire [7:0] coverage_125;
  wire  SaturatingCounter_251_clock;
  wire  SaturatingCounter_251_reset;
  wire  SaturatingCounter_251_io_enable;
  wire  SaturatingCounter_251_io_value;
  wire  _T_1107;
  wire  SaturatingCounter_252_clock;
  wire  SaturatingCounter_252_reset;
  wire  SaturatingCounter_252_io_enable;
  wire  SaturatingCounter_252_io_value;
  wire  _T_1108;
  wire [6:0] _T_1112;
  wire [7:0] coverage_126;
  wire  SaturatingCounter_253_clock;
  wire  SaturatingCounter_253_reset;
  wire  SaturatingCounter_253_io_enable;
  wire  SaturatingCounter_253_io_value;
  wire  _T_1114;
  wire  SaturatingCounter_254_clock;
  wire  SaturatingCounter_254_reset;
  wire  SaturatingCounter_254_io_enable;
  wire  SaturatingCounter_254_io_value;
  wire  _T_1115;
  wire [6:0] _T_1119;
  wire [7:0] coverage_127;
  wire  SaturatingCounter_255_clock;
  wire  SaturatingCounter_255_reset;
  wire  SaturatingCounter_255_io_enable;
  wire  SaturatingCounter_255_io_value;
  wire  _T_1121;
  wire  SaturatingCounter_256_clock;
  wire  SaturatingCounter_256_reset;
  wire  SaturatingCounter_256_io_enable;
  wire  SaturatingCounter_256_io_value;
  wire  _T_1122;
  wire [6:0] _T_1126;
  wire [7:0] coverage_128;
  wire  SaturatingCounter_257_clock;
  wire  SaturatingCounter_257_reset;
  wire  SaturatingCounter_257_io_enable;
  wire  SaturatingCounter_257_io_value;
  wire  _T_1128;
  wire  SaturatingCounter_258_clock;
  wire  SaturatingCounter_258_reset;
  wire  SaturatingCounter_258_io_enable;
  wire  SaturatingCounter_258_io_value;
  wire  _T_1129;
  wire [6:0] _T_1133;
  wire [7:0] coverage_129;
  wire  SaturatingCounter_259_clock;
  wire  SaturatingCounter_259_reset;
  wire  SaturatingCounter_259_io_enable;
  wire  SaturatingCounter_259_io_value;
  wire  _T_1135;
  wire  SaturatingCounter_260_clock;
  wire  SaturatingCounter_260_reset;
  wire  SaturatingCounter_260_io_enable;
  wire  SaturatingCounter_260_io_value;
  wire  _T_1136;
  wire [6:0] _T_1140;
  wire [7:0] coverage_130;
  wire  SaturatingCounter_261_clock;
  wire  SaturatingCounter_261_reset;
  wire  SaturatingCounter_261_io_enable;
  wire  SaturatingCounter_261_io_value;
  wire  _T_1142;
  wire  SaturatingCounter_262_clock;
  wire  SaturatingCounter_262_reset;
  wire  SaturatingCounter_262_io_enable;
  wire  SaturatingCounter_262_io_value;
  wire  _T_1143;
  wire [6:0] _T_1147;
  wire [7:0] coverage_131;
  wire  SaturatingCounter_263_clock;
  wire  SaturatingCounter_263_reset;
  wire  SaturatingCounter_263_io_enable;
  wire  SaturatingCounter_263_io_value;
  wire  _T_1149;
  wire  SaturatingCounter_264_clock;
  wire  SaturatingCounter_264_reset;
  wire  SaturatingCounter_264_io_enable;
  wire  SaturatingCounter_264_io_value;
  wire  _T_1150;
  wire [6:0] _T_1154;
  wire [7:0] coverage_132;
  wire  SaturatingCounter_265_clock;
  wire  SaturatingCounter_265_reset;
  wire  SaturatingCounter_265_io_enable;
  wire  SaturatingCounter_265_io_value;
  wire  _T_1156;
  wire  SaturatingCounter_266_clock;
  wire  SaturatingCounter_266_reset;
  wire  SaturatingCounter_266_io_enable;
  wire  SaturatingCounter_266_io_value;
  wire  _T_1157;
  wire [6:0] _T_1161;
  wire [7:0] coverage_133;
  wire  SaturatingCounter_267_clock;
  wire  SaturatingCounter_267_reset;
  wire  SaturatingCounter_267_io_enable;
  wire  SaturatingCounter_267_io_value;
  wire  _T_1163;
  wire  SaturatingCounter_268_clock;
  wire  SaturatingCounter_268_reset;
  wire  SaturatingCounter_268_io_enable;
  wire  SaturatingCounter_268_io_value;
  wire  _T_1164;
  wire [6:0] _T_1168;
  wire [7:0] coverage_134;
  wire  SaturatingCounter_269_clock;
  wire  SaturatingCounter_269_reset;
  wire  SaturatingCounter_269_io_enable;
  wire  SaturatingCounter_269_io_value;
  wire  _T_1170;
  wire  SaturatingCounter_270_clock;
  wire  SaturatingCounter_270_reset;
  wire  SaturatingCounter_270_io_enable;
  wire  SaturatingCounter_270_io_value;
  wire  _T_1171;
  wire [6:0] _T_1175;
  wire [7:0] coverage_135;
  wire  SaturatingCounter_271_clock;
  wire  SaturatingCounter_271_reset;
  wire  SaturatingCounter_271_io_enable;
  wire  SaturatingCounter_271_io_value;
  wire  _T_1177;
  wire  SaturatingCounter_272_clock;
  wire  SaturatingCounter_272_reset;
  wire  SaturatingCounter_272_io_enable;
  wire  SaturatingCounter_272_io_value;
  wire  _T_1178;
  wire [6:0] _T_1182;
  wire [7:0] coverage_136;
  wire  SaturatingCounter_273_clock;
  wire  SaturatingCounter_273_reset;
  wire  SaturatingCounter_273_io_enable;
  wire  SaturatingCounter_273_io_value;
  wire  _T_1184;
  wire  SaturatingCounter_274_clock;
  wire  SaturatingCounter_274_reset;
  wire  SaturatingCounter_274_io_enable;
  wire  SaturatingCounter_274_io_value;
  wire  _T_1185;
  wire [6:0] _T_1189;
  wire [7:0] coverage_137;
  wire  SaturatingCounter_275_clock;
  wire  SaturatingCounter_275_reset;
  wire  SaturatingCounter_275_io_enable;
  wire  SaturatingCounter_275_io_value;
  wire  _T_1191;
  wire  SaturatingCounter_276_clock;
  wire  SaturatingCounter_276_reset;
  wire  SaturatingCounter_276_io_enable;
  wire  SaturatingCounter_276_io_value;
  wire  _T_1192;
  wire [6:0] _T_1196;
  wire [7:0] coverage_138;
  wire  SaturatingCounter_277_clock;
  wire  SaturatingCounter_277_reset;
  wire  SaturatingCounter_277_io_enable;
  wire  SaturatingCounter_277_io_value;
  wire  _T_1198;
  wire  SaturatingCounter_278_clock;
  wire  SaturatingCounter_278_reset;
  wire  SaturatingCounter_278_io_enable;
  wire  SaturatingCounter_278_io_value;
  wire  _T_1199;
  wire [6:0] _T_1203;
  wire [7:0] coverage_139;
  wire  SaturatingCounter_279_clock;
  wire  SaturatingCounter_279_reset;
  wire  SaturatingCounter_279_io_enable;
  wire  SaturatingCounter_279_io_value;
  wire  _T_1205;
  wire  SaturatingCounter_280_clock;
  wire  SaturatingCounter_280_reset;
  wire  SaturatingCounter_280_io_enable;
  wire  SaturatingCounter_280_io_value;
  wire  _T_1206;
  wire [6:0] _T_1210;
  wire [7:0] coverage_140;
  wire  SaturatingCounter_281_clock;
  wire  SaturatingCounter_281_reset;
  wire  SaturatingCounter_281_io_enable;
  wire  SaturatingCounter_281_io_value;
  wire  _T_1212;
  wire  SaturatingCounter_282_clock;
  wire  SaturatingCounter_282_reset;
  wire  SaturatingCounter_282_io_enable;
  wire  SaturatingCounter_282_io_value;
  wire  _T_1213;
  wire [6:0] _T_1217;
  wire [7:0] coverage_141;
  wire  SaturatingCounter_283_clock;
  wire  SaturatingCounter_283_reset;
  wire  SaturatingCounter_283_io_enable;
  wire  SaturatingCounter_283_io_value;
  wire  _T_1219;
  wire  SaturatingCounter_284_clock;
  wire  SaturatingCounter_284_reset;
  wire  SaturatingCounter_284_io_enable;
  wire  SaturatingCounter_284_io_value;
  wire  _T_1220;
  wire [6:0] _T_1224;
  wire [7:0] coverage_142;
  wire  SaturatingCounter_285_clock;
  wire  SaturatingCounter_285_reset;
  wire  SaturatingCounter_285_io_enable;
  wire  SaturatingCounter_285_io_value;
  wire  _T_1226;
  wire  SaturatingCounter_286_clock;
  wire  SaturatingCounter_286_reset;
  wire  SaturatingCounter_286_io_enable;
  wire  SaturatingCounter_286_io_value;
  wire  _T_1227;
  wire [6:0] _T_1231;
  wire [7:0] coverage_143;
  wire  SaturatingCounter_287_clock;
  wire  SaturatingCounter_287_reset;
  wire  SaturatingCounter_287_io_enable;
  wire  SaturatingCounter_287_io_value;
  wire  _T_1233;
  wire  SaturatingCounter_288_clock;
  wire  SaturatingCounter_288_reset;
  wire  SaturatingCounter_288_io_enable;
  wire  SaturatingCounter_288_io_value;
  wire  _T_1234;
  wire [6:0] _T_1238;
  wire [7:0] coverage_144;
  wire  SaturatingCounter_289_clock;
  wire  SaturatingCounter_289_reset;
  wire  SaturatingCounter_289_io_enable;
  wire  SaturatingCounter_289_io_value;
  wire  _T_1240;
  wire  SaturatingCounter_290_clock;
  wire  SaturatingCounter_290_reset;
  wire  SaturatingCounter_290_io_enable;
  wire  SaturatingCounter_290_io_value;
  wire  _T_1241;
  wire [6:0] _T_1245;
  wire [7:0] coverage_145;
  wire  SaturatingCounter_291_clock;
  wire  SaturatingCounter_291_reset;
  wire  SaturatingCounter_291_io_enable;
  wire  SaturatingCounter_291_io_value;
  wire  _T_1247;
  wire  SaturatingCounter_292_clock;
  wire  SaturatingCounter_292_reset;
  wire  SaturatingCounter_292_io_enable;
  wire  SaturatingCounter_292_io_value;
  wire  _T_1248;
  wire [6:0] _T_1252;
  wire [7:0] coverage_146;
  wire  SaturatingCounter_293_clock;
  wire  SaturatingCounter_293_reset;
  wire  SaturatingCounter_293_io_enable;
  wire  SaturatingCounter_293_io_value;
  wire  _T_1254;
  wire  SaturatingCounter_294_clock;
  wire  SaturatingCounter_294_reset;
  wire  SaturatingCounter_294_io_enable;
  wire  SaturatingCounter_294_io_value;
  wire  _T_1255;
  wire [6:0] _T_1259;
  wire [7:0] coverage_147;
  wire  SaturatingCounter_295_clock;
  wire  SaturatingCounter_295_reset;
  wire  SaturatingCounter_295_io_enable;
  wire  SaturatingCounter_295_io_value;
  wire  _T_1261;
  wire  SaturatingCounter_296_clock;
  wire  SaturatingCounter_296_reset;
  wire  SaturatingCounter_296_io_enable;
  wire  SaturatingCounter_296_io_value;
  wire  _T_1262;
  wire [6:0] _T_1266;
  wire [7:0] coverage_148;
  wire  SaturatingCounter_297_clock;
  wire  SaturatingCounter_297_reset;
  wire  SaturatingCounter_297_io_enable;
  wire  SaturatingCounter_297_io_value;
  wire  _T_1268;
  wire  SaturatingCounter_298_clock;
  wire  SaturatingCounter_298_reset;
  wire  SaturatingCounter_298_io_enable;
  wire  SaturatingCounter_298_io_value;
  wire  _T_1269;
  wire [6:0] _T_1273;
  wire [7:0] coverage_149;
  wire  SaturatingCounter_299_clock;
  wire  SaturatingCounter_299_reset;
  wire  SaturatingCounter_299_io_enable;
  wire  SaturatingCounter_299_io_value;
  wire  _T_1275;
  wire  SaturatingCounter_300_clock;
  wire  SaturatingCounter_300_reset;
  wire  SaturatingCounter_300_io_enable;
  wire  SaturatingCounter_300_io_value;
  wire  _T_1276;
  wire [6:0] _T_1280;
  wire [7:0] coverage_150;
  wire  SaturatingCounter_301_clock;
  wire  SaturatingCounter_301_reset;
  wire  SaturatingCounter_301_io_enable;
  wire  SaturatingCounter_301_io_value;
  wire  _T_1282;
  wire  SaturatingCounter_302_clock;
  wire  SaturatingCounter_302_reset;
  wire  SaturatingCounter_302_io_enable;
  wire  SaturatingCounter_302_io_value;
  wire  _T_1283;
  wire [6:0] _T_1287;
  wire [7:0] coverage_151;
  wire  SaturatingCounter_303_clock;
  wire  SaturatingCounter_303_reset;
  wire  SaturatingCounter_303_io_enable;
  wire  SaturatingCounter_303_io_value;
  wire  _T_1289;
  wire  SaturatingCounter_304_clock;
  wire  SaturatingCounter_304_reset;
  wire  SaturatingCounter_304_io_enable;
  wire  SaturatingCounter_304_io_value;
  wire  _T_1290;
  wire [6:0] _T_1294;
  wire [7:0] coverage_152;
  wire  SaturatingCounter_305_clock;
  wire  SaturatingCounter_305_reset;
  wire  SaturatingCounter_305_io_enable;
  wire  SaturatingCounter_305_io_value;
  wire  _T_1296;
  wire  SaturatingCounter_306_clock;
  wire  SaturatingCounter_306_reset;
  wire  SaturatingCounter_306_io_enable;
  wire  SaturatingCounter_306_io_value;
  wire  _T_1297;
  wire [6:0] _T_1301;
  wire [7:0] coverage_153;
  wire  SaturatingCounter_307_clock;
  wire  SaturatingCounter_307_reset;
  wire  SaturatingCounter_307_io_enable;
  wire  SaturatingCounter_307_io_value;
  wire  _T_1303;
  wire  SaturatingCounter_308_clock;
  wire  SaturatingCounter_308_reset;
  wire  SaturatingCounter_308_io_enable;
  wire  SaturatingCounter_308_io_value;
  wire  _T_1304;
  wire [6:0] _T_1308;
  wire [7:0] coverage_154;
  wire  SaturatingCounter_309_clock;
  wire  SaturatingCounter_309_reset;
  wire  SaturatingCounter_309_io_enable;
  wire  SaturatingCounter_309_io_value;
  wire  _T_1310;
  wire  SaturatingCounter_310_clock;
  wire  SaturatingCounter_310_reset;
  wire  SaturatingCounter_310_io_enable;
  wire  SaturatingCounter_310_io_value;
  wire  _T_1311;
  wire [6:0] _T_1315;
  wire [7:0] coverage_155;
  wire  SaturatingCounter_311_clock;
  wire  SaturatingCounter_311_reset;
  wire  SaturatingCounter_311_io_enable;
  wire  SaturatingCounter_311_io_value;
  wire  _T_1317;
  wire  SaturatingCounter_312_clock;
  wire  SaturatingCounter_312_reset;
  wire  SaturatingCounter_312_io_enable;
  wire  SaturatingCounter_312_io_value;
  wire  _T_1318;
  wire [6:0] _T_1322;
  wire [7:0] coverage_156;
  wire  SaturatingCounter_313_clock;
  wire  SaturatingCounter_313_reset;
  wire  SaturatingCounter_313_io_enable;
  wire  SaturatingCounter_313_io_value;
  wire  _T_1324;
  wire  SaturatingCounter_314_clock;
  wire  SaturatingCounter_314_reset;
  wire  SaturatingCounter_314_io_enable;
  wire  SaturatingCounter_314_io_value;
  wire  _T_1325;
  wire [6:0] _T_1329;
  wire [7:0] coverage_157;
  wire  SaturatingCounter_315_clock;
  wire  SaturatingCounter_315_reset;
  wire  SaturatingCounter_315_io_enable;
  wire  SaturatingCounter_315_io_value;
  wire  _T_1331;
  wire  SaturatingCounter_316_clock;
  wire  SaturatingCounter_316_reset;
  wire  SaturatingCounter_316_io_enable;
  wire  SaturatingCounter_316_io_value;
  wire  _T_1332;
  wire [6:0] _T_1336;
  wire [7:0] coverage_158;
  wire  SaturatingCounter_317_clock;
  wire  SaturatingCounter_317_reset;
  wire  SaturatingCounter_317_io_enable;
  wire  SaturatingCounter_317_io_value;
  wire  _T_1338;
  wire  SaturatingCounter_318_clock;
  wire  SaturatingCounter_318_reset;
  wire  SaturatingCounter_318_io_enable;
  wire  SaturatingCounter_318_io_value;
  wire  _T_1339;
  wire [6:0] _T_1343;
  wire [7:0] coverage_159;
  wire  SaturatingCounter_319_clock;
  wire  SaturatingCounter_319_reset;
  wire  SaturatingCounter_319_io_enable;
  wire  SaturatingCounter_319_io_value;
  wire  _T_1345;
  wire  SaturatingCounter_320_clock;
  wire  SaturatingCounter_320_reset;
  wire  SaturatingCounter_320_io_enable;
  wire  SaturatingCounter_320_io_value;
  wire  _T_1346;
  wire [6:0] _T_1350;
  wire [7:0] coverage_160;
  wire  SaturatingCounter_321_clock;
  wire  SaturatingCounter_321_reset;
  wire  SaturatingCounter_321_io_enable;
  wire  SaturatingCounter_321_io_value;
  wire  _T_1352;
  wire  SaturatingCounter_322_clock;
  wire  SaturatingCounter_322_reset;
  wire  SaturatingCounter_322_io_enable;
  wire  SaturatingCounter_322_io_value;
  wire  _T_1353;
  wire [6:0] _T_1357;
  wire [7:0] coverage_161;
  wire  SaturatingCounter_323_clock;
  wire  SaturatingCounter_323_reset;
  wire  SaturatingCounter_323_io_enable;
  wire  SaturatingCounter_323_io_value;
  wire  _T_1359;
  wire  SaturatingCounter_324_clock;
  wire  SaturatingCounter_324_reset;
  wire  SaturatingCounter_324_io_enable;
  wire  SaturatingCounter_324_io_value;
  wire  _T_1360;
  wire [6:0] _T_1364;
  wire [7:0] coverage_162;
  wire  SaturatingCounter_325_clock;
  wire  SaturatingCounter_325_reset;
  wire  SaturatingCounter_325_io_enable;
  wire  SaturatingCounter_325_io_value;
  wire  _T_1366;
  wire  SaturatingCounter_326_clock;
  wire  SaturatingCounter_326_reset;
  wire  SaturatingCounter_326_io_enable;
  wire  SaturatingCounter_326_io_value;
  wire  _T_1367;
  wire [6:0] _T_1371;
  wire [7:0] coverage_163;
  wire  SaturatingCounter_327_clock;
  wire  SaturatingCounter_327_reset;
  wire  SaturatingCounter_327_io_enable;
  wire  SaturatingCounter_327_io_value;
  wire  _T_1373;
  wire  SaturatingCounter_328_clock;
  wire  SaturatingCounter_328_reset;
  wire  SaturatingCounter_328_io_enable;
  wire  SaturatingCounter_328_io_value;
  wire  _T_1374;
  wire [6:0] _T_1378;
  wire [7:0] coverage_164;
  wire  SaturatingCounter_329_clock;
  wire  SaturatingCounter_329_reset;
  wire  SaturatingCounter_329_io_enable;
  wire  SaturatingCounter_329_io_value;
  wire  _T_1380;
  wire  SaturatingCounter_330_clock;
  wire  SaturatingCounter_330_reset;
  wire  SaturatingCounter_330_io_enable;
  wire  SaturatingCounter_330_io_value;
  wire  _T_1381;
  wire [6:0] _T_1385;
  wire [7:0] coverage_165;
  wire  SaturatingCounter_331_clock;
  wire  SaturatingCounter_331_reset;
  wire  SaturatingCounter_331_io_enable;
  wire  SaturatingCounter_331_io_value;
  wire  _T_1387;
  wire  SaturatingCounter_332_clock;
  wire  SaturatingCounter_332_reset;
  wire  SaturatingCounter_332_io_enable;
  wire  SaturatingCounter_332_io_value;
  wire  _T_1388;
  wire [6:0] _T_1392;
  wire [7:0] coverage_166;
  wire  SaturatingCounter_333_clock;
  wire  SaturatingCounter_333_reset;
  wire  SaturatingCounter_333_io_enable;
  wire  SaturatingCounter_333_io_value;
  wire  _T_1394;
  wire  SaturatingCounter_334_clock;
  wire  SaturatingCounter_334_reset;
  wire  SaturatingCounter_334_io_enable;
  wire  SaturatingCounter_334_io_value;
  wire  _T_1395;
  wire [6:0] _T_1399;
  wire [7:0] coverage_167;
  wire  SaturatingCounter_335_clock;
  wire  SaturatingCounter_335_reset;
  wire  SaturatingCounter_335_io_enable;
  wire  SaturatingCounter_335_io_value;
  wire  _T_1401;
  wire  SaturatingCounter_336_clock;
  wire  SaturatingCounter_336_reset;
  wire  SaturatingCounter_336_io_enable;
  wire  SaturatingCounter_336_io_value;
  wire  _T_1402;
  wire [6:0] _T_1406;
  wire [7:0] coverage_168;
  wire  SaturatingCounter_337_clock;
  wire  SaturatingCounter_337_reset;
  wire  SaturatingCounter_337_io_enable;
  wire  SaturatingCounter_337_io_value;
  wire  _T_1408;
  wire  SaturatingCounter_338_clock;
  wire  SaturatingCounter_338_reset;
  wire  SaturatingCounter_338_io_enable;
  wire  SaturatingCounter_338_io_value;
  wire  _T_1409;
  wire [6:0] _T_1413;
  wire [7:0] coverage_169;
  wire  SaturatingCounter_339_clock;
  wire  SaturatingCounter_339_reset;
  wire  SaturatingCounter_339_io_enable;
  wire  SaturatingCounter_339_io_value;
  wire  _T_1415;
  wire  SaturatingCounter_340_clock;
  wire  SaturatingCounter_340_reset;
  wire  SaturatingCounter_340_io_enable;
  wire  SaturatingCounter_340_io_value;
  wire  _T_1416;
  wire [6:0] _T_1420;
  wire [7:0] coverage_170;
  wire  SaturatingCounter_341_clock;
  wire  SaturatingCounter_341_reset;
  wire  SaturatingCounter_341_io_enable;
  wire  SaturatingCounter_341_io_value;
  wire  _T_1422;
  wire  SaturatingCounter_342_clock;
  wire  SaturatingCounter_342_reset;
  wire  SaturatingCounter_342_io_enable;
  wire  SaturatingCounter_342_io_value;
  wire  _T_1423;
  wire [6:0] _T_1427;
  wire [7:0] coverage_171;
  wire  SaturatingCounter_343_clock;
  wire  SaturatingCounter_343_reset;
  wire  SaturatingCounter_343_io_enable;
  wire  SaturatingCounter_343_io_value;
  wire  _T_1429;
  wire  SaturatingCounter_344_clock;
  wire  SaturatingCounter_344_reset;
  wire  SaturatingCounter_344_io_enable;
  wire  SaturatingCounter_344_io_value;
  wire  _T_1430;
  wire [6:0] _T_1434;
  wire [7:0] coverage_172;
  wire  SaturatingCounter_345_clock;
  wire  SaturatingCounter_345_reset;
  wire  SaturatingCounter_345_io_enable;
  wire  SaturatingCounter_345_io_value;
  wire  _T_1436;
  wire  SaturatingCounter_346_clock;
  wire  SaturatingCounter_346_reset;
  wire  SaturatingCounter_346_io_enable;
  wire  SaturatingCounter_346_io_value;
  wire  _T_1437;
  wire [6:0] _T_1441;
  wire [7:0] coverage_173;
  wire  SaturatingCounter_347_clock;
  wire  SaturatingCounter_347_reset;
  wire  SaturatingCounter_347_io_enable;
  wire  SaturatingCounter_347_io_value;
  wire  _T_1443;
  wire  SaturatingCounter_348_clock;
  wire  SaturatingCounter_348_reset;
  wire  SaturatingCounter_348_io_enable;
  wire  SaturatingCounter_348_io_value;
  wire  _T_1444;
  wire [6:0] _T_1448;
  wire [7:0] coverage_174;
  wire  SaturatingCounter_349_clock;
  wire  SaturatingCounter_349_reset;
  wire  SaturatingCounter_349_io_enable;
  wire  SaturatingCounter_349_io_value;
  wire  _T_1450;
  wire  SaturatingCounter_350_clock;
  wire  SaturatingCounter_350_reset;
  wire  SaturatingCounter_350_io_enable;
  wire  SaturatingCounter_350_io_value;
  wire  _T_1451;
  wire [6:0] _T_1455;
  wire [7:0] coverage_175;
  wire  SaturatingCounter_351_clock;
  wire  SaturatingCounter_351_reset;
  wire  SaturatingCounter_351_io_enable;
  wire  SaturatingCounter_351_io_value;
  wire  _T_1457;
  wire  SaturatingCounter_352_clock;
  wire  SaturatingCounter_352_reset;
  wire  SaturatingCounter_352_io_enable;
  wire  SaturatingCounter_352_io_value;
  wire  _T_1458;
  wire [6:0] _T_1462;
  wire [7:0] coverage_176;
  wire  SaturatingCounter_353_clock;
  wire  SaturatingCounter_353_reset;
  wire  SaturatingCounter_353_io_enable;
  wire  SaturatingCounter_353_io_value;
  wire  _T_1464;
  wire  SaturatingCounter_354_clock;
  wire  SaturatingCounter_354_reset;
  wire  SaturatingCounter_354_io_enable;
  wire  SaturatingCounter_354_io_value;
  wire  _T_1465;
  wire [6:0] _T_1469;
  wire [7:0] coverage_177;
  wire  SaturatingCounter_355_clock;
  wire  SaturatingCounter_355_reset;
  wire  SaturatingCounter_355_io_enable;
  wire  SaturatingCounter_355_io_value;
  wire  _T_1471;
  wire  SaturatingCounter_356_clock;
  wire  SaturatingCounter_356_reset;
  wire  SaturatingCounter_356_io_enable;
  wire  SaturatingCounter_356_io_value;
  wire  _T_1472;
  wire [6:0] _T_1476;
  wire [7:0] coverage_178;
  wire  SaturatingCounter_357_clock;
  wire  SaturatingCounter_357_reset;
  wire  SaturatingCounter_357_io_enable;
  wire  SaturatingCounter_357_io_value;
  wire  _T_1478;
  wire  SaturatingCounter_358_clock;
  wire  SaturatingCounter_358_reset;
  wire  SaturatingCounter_358_io_enable;
  wire  SaturatingCounter_358_io_value;
  wire  _T_1479;
  wire [6:0] _T_1483;
  wire [7:0] coverage_179;
  wire  SaturatingCounter_359_clock;
  wire  SaturatingCounter_359_reset;
  wire  SaturatingCounter_359_io_enable;
  wire  SaturatingCounter_359_io_value;
  wire  _T_1485;
  wire  SaturatingCounter_360_clock;
  wire  SaturatingCounter_360_reset;
  wire  SaturatingCounter_360_io_enable;
  wire  SaturatingCounter_360_io_value;
  wire  _T_1486;
  wire [6:0] _T_1490;
  wire [7:0] coverage_180;
  wire  SaturatingCounter_361_clock;
  wire  SaturatingCounter_361_reset;
  wire  SaturatingCounter_361_io_enable;
  wire  SaturatingCounter_361_io_value;
  wire  _T_1492;
  wire  SaturatingCounter_362_clock;
  wire  SaturatingCounter_362_reset;
  wire  SaturatingCounter_362_io_enable;
  wire  SaturatingCounter_362_io_value;
  wire  _T_1493;
  wire [6:0] _T_1497;
  wire [7:0] coverage_181;
  wire  SaturatingCounter_363_clock;
  wire  SaturatingCounter_363_reset;
  wire  SaturatingCounter_363_io_enable;
  wire  SaturatingCounter_363_io_value;
  wire  _T_1499;
  wire  SaturatingCounter_364_clock;
  wire  SaturatingCounter_364_reset;
  wire  SaturatingCounter_364_io_enable;
  wire  SaturatingCounter_364_io_value;
  wire  _T_1500;
  wire [6:0] _T_1504;
  wire [7:0] coverage_182;
  wire  SaturatingCounter_365_clock;
  wire  SaturatingCounter_365_reset;
  wire  SaturatingCounter_365_io_enable;
  wire  SaturatingCounter_365_io_value;
  wire  _T_1506;
  wire  SaturatingCounter_366_clock;
  wire  SaturatingCounter_366_reset;
  wire  SaturatingCounter_366_io_enable;
  wire  SaturatingCounter_366_io_value;
  wire  _T_1507;
  wire [6:0] _T_1511;
  wire [7:0] coverage_183;
  wire  SaturatingCounter_367_clock;
  wire  SaturatingCounter_367_reset;
  wire  SaturatingCounter_367_io_enable;
  wire  SaturatingCounter_367_io_value;
  wire  _T_1513;
  wire  SaturatingCounter_368_clock;
  wire  SaturatingCounter_368_reset;
  wire  SaturatingCounter_368_io_enable;
  wire  SaturatingCounter_368_io_value;
  wire  _T_1514;
  wire [6:0] _T_1518;
  wire [7:0] coverage_184;
  wire  SaturatingCounter_369_clock;
  wire  SaturatingCounter_369_reset;
  wire  SaturatingCounter_369_io_enable;
  wire  SaturatingCounter_369_io_value;
  wire  _T_1520;
  wire  SaturatingCounter_370_clock;
  wire  SaturatingCounter_370_reset;
  wire  SaturatingCounter_370_io_enable;
  wire  SaturatingCounter_370_io_value;
  wire  _T_1521;
  wire [6:0] _T_1525;
  wire [7:0] coverage_185;
  wire  SaturatingCounter_371_clock;
  wire  SaturatingCounter_371_reset;
  wire  SaturatingCounter_371_io_enable;
  wire  SaturatingCounter_371_io_value;
  wire  _T_1527;
  wire  SaturatingCounter_372_clock;
  wire  SaturatingCounter_372_reset;
  wire  SaturatingCounter_372_io_enable;
  wire  SaturatingCounter_372_io_value;
  wire  _T_1528;
  wire [6:0] _T_1532;
  wire [7:0] coverage_186;
  wire  SaturatingCounter_373_clock;
  wire  SaturatingCounter_373_reset;
  wire  SaturatingCounter_373_io_enable;
  wire  SaturatingCounter_373_io_value;
  wire  _T_1534;
  wire  SaturatingCounter_374_clock;
  wire  SaturatingCounter_374_reset;
  wire  SaturatingCounter_374_io_enable;
  wire  SaturatingCounter_374_io_value;
  wire  _T_1535;
  wire [6:0] _T_1539;
  wire [7:0] coverage_187;
  wire  SaturatingCounter_375_clock;
  wire  SaturatingCounter_375_reset;
  wire  SaturatingCounter_375_io_enable;
  wire  SaturatingCounter_375_io_value;
  wire  _T_1541;
  wire  SaturatingCounter_376_clock;
  wire  SaturatingCounter_376_reset;
  wire  SaturatingCounter_376_io_enable;
  wire  SaturatingCounter_376_io_value;
  wire  _T_1542;
  wire [6:0] _T_1546;
  wire [7:0] coverage_188;
  wire  SaturatingCounter_377_clock;
  wire  SaturatingCounter_377_reset;
  wire  SaturatingCounter_377_io_enable;
  wire  SaturatingCounter_377_io_value;
  wire  _T_1548;
  wire  SaturatingCounter_378_clock;
  wire  SaturatingCounter_378_reset;
  wire  SaturatingCounter_378_io_enable;
  wire  SaturatingCounter_378_io_value;
  wire  _T_1549;
  wire [6:0] _T_1553;
  wire [7:0] coverage_189;
  wire  SaturatingCounter_379_clock;
  wire  SaturatingCounter_379_reset;
  wire  SaturatingCounter_379_io_enable;
  wire  SaturatingCounter_379_io_value;
  wire  _T_1555;
  wire  SaturatingCounter_380_clock;
  wire  SaturatingCounter_380_reset;
  wire  SaturatingCounter_380_io_enable;
  wire  SaturatingCounter_380_io_value;
  wire  _T_1556;
  wire [6:0] _T_1560;
  wire [7:0] coverage_190;
  wire  SaturatingCounter_381_clock;
  wire  SaturatingCounter_381_reset;
  wire  SaturatingCounter_381_io_enable;
  wire  SaturatingCounter_381_io_value;
  wire  _T_1562;
  wire  SaturatingCounter_382_clock;
  wire  SaturatingCounter_382_reset;
  wire  SaturatingCounter_382_io_enable;
  wire  SaturatingCounter_382_io_value;
  wire  _T_1563;
  wire [6:0] _T_1567;
  wire [7:0] coverage_191;
  DUT dut (
    .clock(dut_clock),
    .reset(dut_reset),
    .io_meta_reset(dut_io_meta_reset),
    .io_inputs(dut_io_inputs),
    .io_coverage_0(dut_io_coverage_0),
    .io_coverage_1(dut_io_coverage_1),
    .io_coverage_2(dut_io_coverage_2),
    .io_coverage_3(dut_io_coverage_3),
    .io_coverage_4(dut_io_coverage_4),
    .io_coverage_5(dut_io_coverage_5),
    .io_coverage_6(dut_io_coverage_6),
    .io_coverage_7(dut_io_coverage_7),
    .io_coverage_8(dut_io_coverage_8),
    .io_coverage_9(dut_io_coverage_9),
    .io_coverage_10(dut_io_coverage_10),
    .io_coverage_11(dut_io_coverage_11),
    .io_coverage_12(dut_io_coverage_12),
    .io_coverage_13(dut_io_coverage_13),
    .io_coverage_14(dut_io_coverage_14),
    .io_coverage_15(dut_io_coverage_15),
    .io_coverage_16(dut_io_coverage_16),
    .io_coverage_17(dut_io_coverage_17),
    .io_coverage_18(dut_io_coverage_18),
    .io_coverage_19(dut_io_coverage_19),
    .io_coverage_20(dut_io_coverage_20),
    .io_coverage_21(dut_io_coverage_21),
    .io_coverage_22(dut_io_coverage_22),
    .io_coverage_23(dut_io_coverage_23),
    .io_coverage_24(dut_io_coverage_24),
    .io_coverage_25(dut_io_coverage_25),
    .io_coverage_26(dut_io_coverage_26),
    .io_coverage_27(dut_io_coverage_27),
    .io_coverage_28(dut_io_coverage_28),
    .io_coverage_29(dut_io_coverage_29),
    .io_coverage_30(dut_io_coverage_30),
    .io_coverage_31(dut_io_coverage_31),
    .io_coverage_32(dut_io_coverage_32),
    .io_coverage_33(dut_io_coverage_33),
    .io_coverage_34(dut_io_coverage_34),
    .io_coverage_35(dut_io_coverage_35),
    .io_coverage_36(dut_io_coverage_36),
    .io_coverage_37(dut_io_coverage_37),
    .io_coverage_38(dut_io_coverage_38),
    .io_coverage_39(dut_io_coverage_39),
    .io_coverage_40(dut_io_coverage_40),
    .io_coverage_41(dut_io_coverage_41),
    .io_coverage_42(dut_io_coverage_42),
    .io_coverage_43(dut_io_coverage_43),
    .io_coverage_44(dut_io_coverage_44),
    .io_coverage_45(dut_io_coverage_45),
    .io_coverage_46(dut_io_coverage_46),
    .io_coverage_47(dut_io_coverage_47),
    .io_coverage_48(dut_io_coverage_48),
    .io_coverage_49(dut_io_coverage_49),
    .io_coverage_50(dut_io_coverage_50),
    .io_coverage_51(dut_io_coverage_51),
    .io_coverage_52(dut_io_coverage_52),
    .io_coverage_53(dut_io_coverage_53),
    .io_coverage_54(dut_io_coverage_54),
    .io_coverage_55(dut_io_coverage_55),
    .io_coverage_56(dut_io_coverage_56),
    .io_coverage_57(dut_io_coverage_57),
    .io_coverage_58(dut_io_coverage_58),
    .io_coverage_59(dut_io_coverage_59),
    .io_coverage_60(dut_io_coverage_60),
    .io_coverage_61(dut_io_coverage_61),
    .io_coverage_62(dut_io_coverage_62),
    .io_coverage_63(dut_io_coverage_63),
    .io_coverage_64(dut_io_coverage_64),
    .io_coverage_65(dut_io_coverage_65),
    .io_coverage_66(dut_io_coverage_66),
    .io_coverage_67(dut_io_coverage_67),
    .io_coverage_68(dut_io_coverage_68),
    .io_coverage_69(dut_io_coverage_69),
    .io_coverage_70(dut_io_coverage_70),
    .io_coverage_71(dut_io_coverage_71),
    .io_coverage_72(dut_io_coverage_72),
    .io_coverage_73(dut_io_coverage_73),
    .io_coverage_74(dut_io_coverage_74),
    .io_coverage_75(dut_io_coverage_75),
    .io_coverage_76(dut_io_coverage_76),
    .io_coverage_77(dut_io_coverage_77),
    .io_coverage_78(dut_io_coverage_78),
    .io_coverage_79(dut_io_coverage_79),
    .io_coverage_80(dut_io_coverage_80),
    .io_coverage_81(dut_io_coverage_81),
    .io_coverage_82(dut_io_coverage_82),
    .io_coverage_83(dut_io_coverage_83),
    .io_coverage_84(dut_io_coverage_84),
    .io_coverage_85(dut_io_coverage_85),
    .io_coverage_86(dut_io_coverage_86),
    .io_coverage_87(dut_io_coverage_87),
    .io_coverage_88(dut_io_coverage_88),
    .io_coverage_89(dut_io_coverage_89),
    .io_coverage_90(dut_io_coverage_90),
    .io_coverage_91(dut_io_coverage_91),
    .io_coverage_92(dut_io_coverage_92),
    .io_coverage_93(dut_io_coverage_93),
    .io_coverage_94(dut_io_coverage_94),
    .io_coverage_95(dut_io_coverage_95),
    .io_coverage_96(dut_io_coverage_96),
    .io_coverage_97(dut_io_coverage_97),
    .io_coverage_98(dut_io_coverage_98),
    .io_coverage_99(dut_io_coverage_99),
    .io_coverage_100(dut_io_coverage_100),
    .io_coverage_101(dut_io_coverage_101),
    .io_coverage_102(dut_io_coverage_102),
    .io_coverage_103(dut_io_coverage_103),
    .io_coverage_104(dut_io_coverage_104),
    .io_coverage_105(dut_io_coverage_105),
    .io_coverage_106(dut_io_coverage_106),
    .io_coverage_107(dut_io_coverage_107),
    .io_coverage_108(dut_io_coverage_108),
    .io_coverage_109(dut_io_coverage_109),
    .io_coverage_110(dut_io_coverage_110),
    .io_coverage_111(dut_io_coverage_111),
    .io_coverage_112(dut_io_coverage_112),
    .io_coverage_113(dut_io_coverage_113),
    .io_coverage_114(dut_io_coverage_114),
    .io_coverage_115(dut_io_coverage_115),
    .io_coverage_116(dut_io_coverage_116),
    .io_coverage_117(dut_io_coverage_117),
    .io_coverage_118(dut_io_coverage_118),
    .io_coverage_119(dut_io_coverage_119),
    .io_coverage_120(dut_io_coverage_120),
    .io_coverage_121(dut_io_coverage_121),
    .io_coverage_122(dut_io_coverage_122),
    .io_coverage_123(dut_io_coverage_123),
    .io_coverage_124(dut_io_coverage_124),
    .io_coverage_125(dut_io_coverage_125),
    .io_coverage_126(dut_io_coverage_126),
    .io_coverage_127(dut_io_coverage_127),
    .io_coverage_128(dut_io_coverage_128),
    .io_coverage_129(dut_io_coverage_129),
    .io_coverage_130(dut_io_coverage_130),
    .io_coverage_131(dut_io_coverage_131),
    .io_coverage_132(dut_io_coverage_132),
    .io_coverage_133(dut_io_coverage_133),
    .io_coverage_134(dut_io_coverage_134),
    .io_coverage_135(dut_io_coverage_135),
    .io_coverage_136(dut_io_coverage_136),
    .io_coverage_137(dut_io_coverage_137),
    .io_coverage_138(dut_io_coverage_138),
    .io_coverage_139(dut_io_coverage_139),
    .io_coverage_140(dut_io_coverage_140),
    .io_coverage_141(dut_io_coverage_141),
    .io_coverage_142(dut_io_coverage_142),
    .io_coverage_143(dut_io_coverage_143),
    .io_coverage_144(dut_io_coverage_144),
    .io_coverage_145(dut_io_coverage_145),
    .io_coverage_146(dut_io_coverage_146),
    .io_coverage_147(dut_io_coverage_147),
    .io_coverage_148(dut_io_coverage_148),
    .io_coverage_149(dut_io_coverage_149),
    .io_coverage_150(dut_io_coverage_150),
    .io_coverage_151(dut_io_coverage_151),
    .io_coverage_152(dut_io_coverage_152),
    .io_coverage_153(dut_io_coverage_153),
    .io_coverage_154(dut_io_coverage_154),
    .io_coverage_155(dut_io_coverage_155),
    .io_coverage_156(dut_io_coverage_156),
    .io_coverage_157(dut_io_coverage_157),
    .io_coverage_158(dut_io_coverage_158),
    .io_coverage_159(dut_io_coverage_159),
    .io_coverage_160(dut_io_coverage_160),
    .io_coverage_161(dut_io_coverage_161),
    .io_coverage_162(dut_io_coverage_162),
    .io_coverage_163(dut_io_coverage_163),
    .io_coverage_164(dut_io_coverage_164),
    .io_coverage_165(dut_io_coverage_165),
    .io_coverage_166(dut_io_coverage_166),
    .io_coverage_167(dut_io_coverage_167),
    .io_coverage_168(dut_io_coverage_168),
    .io_coverage_169(dut_io_coverage_169),
    .io_coverage_170(dut_io_coverage_170),
    .io_coverage_171(dut_io_coverage_171),
    .io_coverage_172(dut_io_coverage_172),
    .io_coverage_173(dut_io_coverage_173),
    .io_coverage_174(dut_io_coverage_174),
    .io_coverage_175(dut_io_coverage_175),
    .io_coverage_176(dut_io_coverage_176),
    .io_coverage_177(dut_io_coverage_177),
    .io_coverage_178(dut_io_coverage_178),
    .io_coverage_179(dut_io_coverage_179),
    .io_coverage_180(dut_io_coverage_180),
    .io_coverage_181(dut_io_coverage_181),
    .io_coverage_182(dut_io_coverage_182),
    .io_coverage_183(dut_io_coverage_183),
    .io_coverage_184(dut_io_coverage_184),
    .io_coverage_185(dut_io_coverage_185),
    .io_coverage_186(dut_io_coverage_186),
    .io_coverage_187(dut_io_coverage_187),
    .io_coverage_188(dut_io_coverage_188),
    .io_coverage_189(dut_io_coverage_189),
    .io_coverage_190(dut_io_coverage_190),
    .io_coverage_191(dut_io_coverage_191)
  );
  SaturatingCounter SaturatingCounter (
    .clock(SaturatingCounter_clock),
    .reset(SaturatingCounter_reset),
    .io_enable(SaturatingCounter_io_enable),
    .io_value(SaturatingCounter_io_value)
  );
  SaturatingCounter SaturatingCounter_1 (
    .clock(SaturatingCounter_1_clock),
    .reset(SaturatingCounter_1_reset),
    .io_enable(SaturatingCounter_1_io_enable),
    .io_value(SaturatingCounter_1_io_value)
  );
  SaturatingCounter SaturatingCounter_2 (
    .clock(SaturatingCounter_2_clock),
    .reset(SaturatingCounter_2_reset),
    .io_enable(SaturatingCounter_2_io_enable),
    .io_value(SaturatingCounter_2_io_value)
  );
  SaturatingCounter SaturatingCounter_3 (
    .clock(SaturatingCounter_3_clock),
    .reset(SaturatingCounter_3_reset),
    .io_enable(SaturatingCounter_3_io_enable),
    .io_value(SaturatingCounter_3_io_value)
  );
  SaturatingCounter SaturatingCounter_4 (
    .clock(SaturatingCounter_4_clock),
    .reset(SaturatingCounter_4_reset),
    .io_enable(SaturatingCounter_4_io_enable),
    .io_value(SaturatingCounter_4_io_value)
  );
  SaturatingCounter SaturatingCounter_5 (
    .clock(SaturatingCounter_5_clock),
    .reset(SaturatingCounter_5_reset),
    .io_enable(SaturatingCounter_5_io_enable),
    .io_value(SaturatingCounter_5_io_value)
  );
  SaturatingCounter SaturatingCounter_6 (
    .clock(SaturatingCounter_6_clock),
    .reset(SaturatingCounter_6_reset),
    .io_enable(SaturatingCounter_6_io_enable),
    .io_value(SaturatingCounter_6_io_value)
  );
  SaturatingCounter SaturatingCounter_7 (
    .clock(SaturatingCounter_7_clock),
    .reset(SaturatingCounter_7_reset),
    .io_enable(SaturatingCounter_7_io_enable),
    .io_value(SaturatingCounter_7_io_value)
  );
  SaturatingCounter SaturatingCounter_8 (
    .clock(SaturatingCounter_8_clock),
    .reset(SaturatingCounter_8_reset),
    .io_enable(SaturatingCounter_8_io_enable),
    .io_value(SaturatingCounter_8_io_value)
  );
  SaturatingCounter SaturatingCounter_9 (
    .clock(SaturatingCounter_9_clock),
    .reset(SaturatingCounter_9_reset),
    .io_enable(SaturatingCounter_9_io_enable),
    .io_value(SaturatingCounter_9_io_value)
  );
  SaturatingCounter SaturatingCounter_10 (
    .clock(SaturatingCounter_10_clock),
    .reset(SaturatingCounter_10_reset),
    .io_enable(SaturatingCounter_10_io_enable),
    .io_value(SaturatingCounter_10_io_value)
  );
  SaturatingCounter SaturatingCounter_11 (
    .clock(SaturatingCounter_11_clock),
    .reset(SaturatingCounter_11_reset),
    .io_enable(SaturatingCounter_11_io_enable),
    .io_value(SaturatingCounter_11_io_value)
  );
  SaturatingCounter SaturatingCounter_12 (
    .clock(SaturatingCounter_12_clock),
    .reset(SaturatingCounter_12_reset),
    .io_enable(SaturatingCounter_12_io_enable),
    .io_value(SaturatingCounter_12_io_value)
  );
  SaturatingCounter SaturatingCounter_13 (
    .clock(SaturatingCounter_13_clock),
    .reset(SaturatingCounter_13_reset),
    .io_enable(SaturatingCounter_13_io_enable),
    .io_value(SaturatingCounter_13_io_value)
  );
  SaturatingCounter SaturatingCounter_14 (
    .clock(SaturatingCounter_14_clock),
    .reset(SaturatingCounter_14_reset),
    .io_enable(SaturatingCounter_14_io_enable),
    .io_value(SaturatingCounter_14_io_value)
  );
  SaturatingCounter SaturatingCounter_15 (
    .clock(SaturatingCounter_15_clock),
    .reset(SaturatingCounter_15_reset),
    .io_enable(SaturatingCounter_15_io_enable),
    .io_value(SaturatingCounter_15_io_value)
  );
  SaturatingCounter SaturatingCounter_16 (
    .clock(SaturatingCounter_16_clock),
    .reset(SaturatingCounter_16_reset),
    .io_enable(SaturatingCounter_16_io_enable),
    .io_value(SaturatingCounter_16_io_value)
  );
  SaturatingCounter SaturatingCounter_17 (
    .clock(SaturatingCounter_17_clock),
    .reset(SaturatingCounter_17_reset),
    .io_enable(SaturatingCounter_17_io_enable),
    .io_value(SaturatingCounter_17_io_value)
  );
  SaturatingCounter SaturatingCounter_18 (
    .clock(SaturatingCounter_18_clock),
    .reset(SaturatingCounter_18_reset),
    .io_enable(SaturatingCounter_18_io_enable),
    .io_value(SaturatingCounter_18_io_value)
  );
  SaturatingCounter SaturatingCounter_19 (
    .clock(SaturatingCounter_19_clock),
    .reset(SaturatingCounter_19_reset),
    .io_enable(SaturatingCounter_19_io_enable),
    .io_value(SaturatingCounter_19_io_value)
  );
  SaturatingCounter SaturatingCounter_20 (
    .clock(SaturatingCounter_20_clock),
    .reset(SaturatingCounter_20_reset),
    .io_enable(SaturatingCounter_20_io_enable),
    .io_value(SaturatingCounter_20_io_value)
  );
  SaturatingCounter SaturatingCounter_21 (
    .clock(SaturatingCounter_21_clock),
    .reset(SaturatingCounter_21_reset),
    .io_enable(SaturatingCounter_21_io_enable),
    .io_value(SaturatingCounter_21_io_value)
  );
  SaturatingCounter SaturatingCounter_22 (
    .clock(SaturatingCounter_22_clock),
    .reset(SaturatingCounter_22_reset),
    .io_enable(SaturatingCounter_22_io_enable),
    .io_value(SaturatingCounter_22_io_value)
  );
  SaturatingCounter SaturatingCounter_23 (
    .clock(SaturatingCounter_23_clock),
    .reset(SaturatingCounter_23_reset),
    .io_enable(SaturatingCounter_23_io_enable),
    .io_value(SaturatingCounter_23_io_value)
  );
  SaturatingCounter SaturatingCounter_24 (
    .clock(SaturatingCounter_24_clock),
    .reset(SaturatingCounter_24_reset),
    .io_enable(SaturatingCounter_24_io_enable),
    .io_value(SaturatingCounter_24_io_value)
  );
  SaturatingCounter SaturatingCounter_25 (
    .clock(SaturatingCounter_25_clock),
    .reset(SaturatingCounter_25_reset),
    .io_enable(SaturatingCounter_25_io_enable),
    .io_value(SaturatingCounter_25_io_value)
  );
  SaturatingCounter SaturatingCounter_26 (
    .clock(SaturatingCounter_26_clock),
    .reset(SaturatingCounter_26_reset),
    .io_enable(SaturatingCounter_26_io_enable),
    .io_value(SaturatingCounter_26_io_value)
  );
  SaturatingCounter SaturatingCounter_27 (
    .clock(SaturatingCounter_27_clock),
    .reset(SaturatingCounter_27_reset),
    .io_enable(SaturatingCounter_27_io_enable),
    .io_value(SaturatingCounter_27_io_value)
  );
  SaturatingCounter SaturatingCounter_28 (
    .clock(SaturatingCounter_28_clock),
    .reset(SaturatingCounter_28_reset),
    .io_enable(SaturatingCounter_28_io_enable),
    .io_value(SaturatingCounter_28_io_value)
  );
  SaturatingCounter SaturatingCounter_29 (
    .clock(SaturatingCounter_29_clock),
    .reset(SaturatingCounter_29_reset),
    .io_enable(SaturatingCounter_29_io_enable),
    .io_value(SaturatingCounter_29_io_value)
  );
  SaturatingCounter SaturatingCounter_30 (
    .clock(SaturatingCounter_30_clock),
    .reset(SaturatingCounter_30_reset),
    .io_enable(SaturatingCounter_30_io_enable),
    .io_value(SaturatingCounter_30_io_value)
  );
  SaturatingCounter SaturatingCounter_31 (
    .clock(SaturatingCounter_31_clock),
    .reset(SaturatingCounter_31_reset),
    .io_enable(SaturatingCounter_31_io_enable),
    .io_value(SaturatingCounter_31_io_value)
  );
  SaturatingCounter SaturatingCounter_32 (
    .clock(SaturatingCounter_32_clock),
    .reset(SaturatingCounter_32_reset),
    .io_enable(SaturatingCounter_32_io_enable),
    .io_value(SaturatingCounter_32_io_value)
  );
  SaturatingCounter SaturatingCounter_33 (
    .clock(SaturatingCounter_33_clock),
    .reset(SaturatingCounter_33_reset),
    .io_enable(SaturatingCounter_33_io_enable),
    .io_value(SaturatingCounter_33_io_value)
  );
  SaturatingCounter SaturatingCounter_34 (
    .clock(SaturatingCounter_34_clock),
    .reset(SaturatingCounter_34_reset),
    .io_enable(SaturatingCounter_34_io_enable),
    .io_value(SaturatingCounter_34_io_value)
  );
  SaturatingCounter SaturatingCounter_35 (
    .clock(SaturatingCounter_35_clock),
    .reset(SaturatingCounter_35_reset),
    .io_enable(SaturatingCounter_35_io_enable),
    .io_value(SaturatingCounter_35_io_value)
  );
  SaturatingCounter SaturatingCounter_36 (
    .clock(SaturatingCounter_36_clock),
    .reset(SaturatingCounter_36_reset),
    .io_enable(SaturatingCounter_36_io_enable),
    .io_value(SaturatingCounter_36_io_value)
  );
  SaturatingCounter SaturatingCounter_37 (
    .clock(SaturatingCounter_37_clock),
    .reset(SaturatingCounter_37_reset),
    .io_enable(SaturatingCounter_37_io_enable),
    .io_value(SaturatingCounter_37_io_value)
  );
  SaturatingCounter SaturatingCounter_38 (
    .clock(SaturatingCounter_38_clock),
    .reset(SaturatingCounter_38_reset),
    .io_enable(SaturatingCounter_38_io_enable),
    .io_value(SaturatingCounter_38_io_value)
  );
  SaturatingCounter SaturatingCounter_39 (
    .clock(SaturatingCounter_39_clock),
    .reset(SaturatingCounter_39_reset),
    .io_enable(SaturatingCounter_39_io_enable),
    .io_value(SaturatingCounter_39_io_value)
  );
  SaturatingCounter SaturatingCounter_40 (
    .clock(SaturatingCounter_40_clock),
    .reset(SaturatingCounter_40_reset),
    .io_enable(SaturatingCounter_40_io_enable),
    .io_value(SaturatingCounter_40_io_value)
  );
  SaturatingCounter SaturatingCounter_41 (
    .clock(SaturatingCounter_41_clock),
    .reset(SaturatingCounter_41_reset),
    .io_enable(SaturatingCounter_41_io_enable),
    .io_value(SaturatingCounter_41_io_value)
  );
  SaturatingCounter SaturatingCounter_42 (
    .clock(SaturatingCounter_42_clock),
    .reset(SaturatingCounter_42_reset),
    .io_enable(SaturatingCounter_42_io_enable),
    .io_value(SaturatingCounter_42_io_value)
  );
  SaturatingCounter SaturatingCounter_43 (
    .clock(SaturatingCounter_43_clock),
    .reset(SaturatingCounter_43_reset),
    .io_enable(SaturatingCounter_43_io_enable),
    .io_value(SaturatingCounter_43_io_value)
  );
  SaturatingCounter SaturatingCounter_44 (
    .clock(SaturatingCounter_44_clock),
    .reset(SaturatingCounter_44_reset),
    .io_enable(SaturatingCounter_44_io_enable),
    .io_value(SaturatingCounter_44_io_value)
  );
  SaturatingCounter SaturatingCounter_45 (
    .clock(SaturatingCounter_45_clock),
    .reset(SaturatingCounter_45_reset),
    .io_enable(SaturatingCounter_45_io_enable),
    .io_value(SaturatingCounter_45_io_value)
  );
  SaturatingCounter SaturatingCounter_46 (
    .clock(SaturatingCounter_46_clock),
    .reset(SaturatingCounter_46_reset),
    .io_enable(SaturatingCounter_46_io_enable),
    .io_value(SaturatingCounter_46_io_value)
  );
  SaturatingCounter SaturatingCounter_47 (
    .clock(SaturatingCounter_47_clock),
    .reset(SaturatingCounter_47_reset),
    .io_enable(SaturatingCounter_47_io_enable),
    .io_value(SaturatingCounter_47_io_value)
  );
  SaturatingCounter SaturatingCounter_48 (
    .clock(SaturatingCounter_48_clock),
    .reset(SaturatingCounter_48_reset),
    .io_enable(SaturatingCounter_48_io_enable),
    .io_value(SaturatingCounter_48_io_value)
  );
  SaturatingCounter SaturatingCounter_49 (
    .clock(SaturatingCounter_49_clock),
    .reset(SaturatingCounter_49_reset),
    .io_enable(SaturatingCounter_49_io_enable),
    .io_value(SaturatingCounter_49_io_value)
  );
  SaturatingCounter SaturatingCounter_50 (
    .clock(SaturatingCounter_50_clock),
    .reset(SaturatingCounter_50_reset),
    .io_enable(SaturatingCounter_50_io_enable),
    .io_value(SaturatingCounter_50_io_value)
  );
  SaturatingCounter SaturatingCounter_51 (
    .clock(SaturatingCounter_51_clock),
    .reset(SaturatingCounter_51_reset),
    .io_enable(SaturatingCounter_51_io_enable),
    .io_value(SaturatingCounter_51_io_value)
  );
  SaturatingCounter SaturatingCounter_52 (
    .clock(SaturatingCounter_52_clock),
    .reset(SaturatingCounter_52_reset),
    .io_enable(SaturatingCounter_52_io_enable),
    .io_value(SaturatingCounter_52_io_value)
  );
  SaturatingCounter SaturatingCounter_53 (
    .clock(SaturatingCounter_53_clock),
    .reset(SaturatingCounter_53_reset),
    .io_enable(SaturatingCounter_53_io_enable),
    .io_value(SaturatingCounter_53_io_value)
  );
  SaturatingCounter SaturatingCounter_54 (
    .clock(SaturatingCounter_54_clock),
    .reset(SaturatingCounter_54_reset),
    .io_enable(SaturatingCounter_54_io_enable),
    .io_value(SaturatingCounter_54_io_value)
  );
  SaturatingCounter SaturatingCounter_55 (
    .clock(SaturatingCounter_55_clock),
    .reset(SaturatingCounter_55_reset),
    .io_enable(SaturatingCounter_55_io_enable),
    .io_value(SaturatingCounter_55_io_value)
  );
  SaturatingCounter SaturatingCounter_56 (
    .clock(SaturatingCounter_56_clock),
    .reset(SaturatingCounter_56_reset),
    .io_enable(SaturatingCounter_56_io_enable),
    .io_value(SaturatingCounter_56_io_value)
  );
  SaturatingCounter SaturatingCounter_57 (
    .clock(SaturatingCounter_57_clock),
    .reset(SaturatingCounter_57_reset),
    .io_enable(SaturatingCounter_57_io_enable),
    .io_value(SaturatingCounter_57_io_value)
  );
  SaturatingCounter SaturatingCounter_58 (
    .clock(SaturatingCounter_58_clock),
    .reset(SaturatingCounter_58_reset),
    .io_enable(SaturatingCounter_58_io_enable),
    .io_value(SaturatingCounter_58_io_value)
  );
  SaturatingCounter SaturatingCounter_59 (
    .clock(SaturatingCounter_59_clock),
    .reset(SaturatingCounter_59_reset),
    .io_enable(SaturatingCounter_59_io_enable),
    .io_value(SaturatingCounter_59_io_value)
  );
  SaturatingCounter SaturatingCounter_60 (
    .clock(SaturatingCounter_60_clock),
    .reset(SaturatingCounter_60_reset),
    .io_enable(SaturatingCounter_60_io_enable),
    .io_value(SaturatingCounter_60_io_value)
  );
  SaturatingCounter SaturatingCounter_61 (
    .clock(SaturatingCounter_61_clock),
    .reset(SaturatingCounter_61_reset),
    .io_enable(SaturatingCounter_61_io_enable),
    .io_value(SaturatingCounter_61_io_value)
  );
  SaturatingCounter SaturatingCounter_62 (
    .clock(SaturatingCounter_62_clock),
    .reset(SaturatingCounter_62_reset),
    .io_enable(SaturatingCounter_62_io_enable),
    .io_value(SaturatingCounter_62_io_value)
  );
  SaturatingCounter SaturatingCounter_63 (
    .clock(SaturatingCounter_63_clock),
    .reset(SaturatingCounter_63_reset),
    .io_enable(SaturatingCounter_63_io_enable),
    .io_value(SaturatingCounter_63_io_value)
  );
  SaturatingCounter SaturatingCounter_64 (
    .clock(SaturatingCounter_64_clock),
    .reset(SaturatingCounter_64_reset),
    .io_enable(SaturatingCounter_64_io_enable),
    .io_value(SaturatingCounter_64_io_value)
  );
  SaturatingCounter SaturatingCounter_65 (
    .clock(SaturatingCounter_65_clock),
    .reset(SaturatingCounter_65_reset),
    .io_enable(SaturatingCounter_65_io_enable),
    .io_value(SaturatingCounter_65_io_value)
  );
  SaturatingCounter SaturatingCounter_66 (
    .clock(SaturatingCounter_66_clock),
    .reset(SaturatingCounter_66_reset),
    .io_enable(SaturatingCounter_66_io_enable),
    .io_value(SaturatingCounter_66_io_value)
  );
  SaturatingCounter SaturatingCounter_67 (
    .clock(SaturatingCounter_67_clock),
    .reset(SaturatingCounter_67_reset),
    .io_enable(SaturatingCounter_67_io_enable),
    .io_value(SaturatingCounter_67_io_value)
  );
  SaturatingCounter SaturatingCounter_68 (
    .clock(SaturatingCounter_68_clock),
    .reset(SaturatingCounter_68_reset),
    .io_enable(SaturatingCounter_68_io_enable),
    .io_value(SaturatingCounter_68_io_value)
  );
  SaturatingCounter SaturatingCounter_69 (
    .clock(SaturatingCounter_69_clock),
    .reset(SaturatingCounter_69_reset),
    .io_enable(SaturatingCounter_69_io_enable),
    .io_value(SaturatingCounter_69_io_value)
  );
  SaturatingCounter SaturatingCounter_70 (
    .clock(SaturatingCounter_70_clock),
    .reset(SaturatingCounter_70_reset),
    .io_enable(SaturatingCounter_70_io_enable),
    .io_value(SaturatingCounter_70_io_value)
  );
  SaturatingCounter SaturatingCounter_71 (
    .clock(SaturatingCounter_71_clock),
    .reset(SaturatingCounter_71_reset),
    .io_enable(SaturatingCounter_71_io_enable),
    .io_value(SaturatingCounter_71_io_value)
  );
  SaturatingCounter SaturatingCounter_72 (
    .clock(SaturatingCounter_72_clock),
    .reset(SaturatingCounter_72_reset),
    .io_enable(SaturatingCounter_72_io_enable),
    .io_value(SaturatingCounter_72_io_value)
  );
  SaturatingCounter SaturatingCounter_73 (
    .clock(SaturatingCounter_73_clock),
    .reset(SaturatingCounter_73_reset),
    .io_enable(SaturatingCounter_73_io_enable),
    .io_value(SaturatingCounter_73_io_value)
  );
  SaturatingCounter SaturatingCounter_74 (
    .clock(SaturatingCounter_74_clock),
    .reset(SaturatingCounter_74_reset),
    .io_enable(SaturatingCounter_74_io_enable),
    .io_value(SaturatingCounter_74_io_value)
  );
  SaturatingCounter SaturatingCounter_75 (
    .clock(SaturatingCounter_75_clock),
    .reset(SaturatingCounter_75_reset),
    .io_enable(SaturatingCounter_75_io_enable),
    .io_value(SaturatingCounter_75_io_value)
  );
  SaturatingCounter SaturatingCounter_76 (
    .clock(SaturatingCounter_76_clock),
    .reset(SaturatingCounter_76_reset),
    .io_enable(SaturatingCounter_76_io_enable),
    .io_value(SaturatingCounter_76_io_value)
  );
  SaturatingCounter SaturatingCounter_77 (
    .clock(SaturatingCounter_77_clock),
    .reset(SaturatingCounter_77_reset),
    .io_enable(SaturatingCounter_77_io_enable),
    .io_value(SaturatingCounter_77_io_value)
  );
  SaturatingCounter SaturatingCounter_78 (
    .clock(SaturatingCounter_78_clock),
    .reset(SaturatingCounter_78_reset),
    .io_enable(SaturatingCounter_78_io_enable),
    .io_value(SaturatingCounter_78_io_value)
  );
  SaturatingCounter SaturatingCounter_79 (
    .clock(SaturatingCounter_79_clock),
    .reset(SaturatingCounter_79_reset),
    .io_enable(SaturatingCounter_79_io_enable),
    .io_value(SaturatingCounter_79_io_value)
  );
  SaturatingCounter SaturatingCounter_80 (
    .clock(SaturatingCounter_80_clock),
    .reset(SaturatingCounter_80_reset),
    .io_enable(SaturatingCounter_80_io_enable),
    .io_value(SaturatingCounter_80_io_value)
  );
  SaturatingCounter SaturatingCounter_81 (
    .clock(SaturatingCounter_81_clock),
    .reset(SaturatingCounter_81_reset),
    .io_enable(SaturatingCounter_81_io_enable),
    .io_value(SaturatingCounter_81_io_value)
  );
  SaturatingCounter SaturatingCounter_82 (
    .clock(SaturatingCounter_82_clock),
    .reset(SaturatingCounter_82_reset),
    .io_enable(SaturatingCounter_82_io_enable),
    .io_value(SaturatingCounter_82_io_value)
  );
  SaturatingCounter SaturatingCounter_83 (
    .clock(SaturatingCounter_83_clock),
    .reset(SaturatingCounter_83_reset),
    .io_enable(SaturatingCounter_83_io_enable),
    .io_value(SaturatingCounter_83_io_value)
  );
  SaturatingCounter SaturatingCounter_84 (
    .clock(SaturatingCounter_84_clock),
    .reset(SaturatingCounter_84_reset),
    .io_enable(SaturatingCounter_84_io_enable),
    .io_value(SaturatingCounter_84_io_value)
  );
  SaturatingCounter SaturatingCounter_85 (
    .clock(SaturatingCounter_85_clock),
    .reset(SaturatingCounter_85_reset),
    .io_enable(SaturatingCounter_85_io_enable),
    .io_value(SaturatingCounter_85_io_value)
  );
  SaturatingCounter SaturatingCounter_86 (
    .clock(SaturatingCounter_86_clock),
    .reset(SaturatingCounter_86_reset),
    .io_enable(SaturatingCounter_86_io_enable),
    .io_value(SaturatingCounter_86_io_value)
  );
  SaturatingCounter SaturatingCounter_87 (
    .clock(SaturatingCounter_87_clock),
    .reset(SaturatingCounter_87_reset),
    .io_enable(SaturatingCounter_87_io_enable),
    .io_value(SaturatingCounter_87_io_value)
  );
  SaturatingCounter SaturatingCounter_88 (
    .clock(SaturatingCounter_88_clock),
    .reset(SaturatingCounter_88_reset),
    .io_enable(SaturatingCounter_88_io_enable),
    .io_value(SaturatingCounter_88_io_value)
  );
  SaturatingCounter SaturatingCounter_89 (
    .clock(SaturatingCounter_89_clock),
    .reset(SaturatingCounter_89_reset),
    .io_enable(SaturatingCounter_89_io_enable),
    .io_value(SaturatingCounter_89_io_value)
  );
  SaturatingCounter SaturatingCounter_90 (
    .clock(SaturatingCounter_90_clock),
    .reset(SaturatingCounter_90_reset),
    .io_enable(SaturatingCounter_90_io_enable),
    .io_value(SaturatingCounter_90_io_value)
  );
  SaturatingCounter SaturatingCounter_91 (
    .clock(SaturatingCounter_91_clock),
    .reset(SaturatingCounter_91_reset),
    .io_enable(SaturatingCounter_91_io_enable),
    .io_value(SaturatingCounter_91_io_value)
  );
  SaturatingCounter SaturatingCounter_92 (
    .clock(SaturatingCounter_92_clock),
    .reset(SaturatingCounter_92_reset),
    .io_enable(SaturatingCounter_92_io_enable),
    .io_value(SaturatingCounter_92_io_value)
  );
  SaturatingCounter SaturatingCounter_93 (
    .clock(SaturatingCounter_93_clock),
    .reset(SaturatingCounter_93_reset),
    .io_enable(SaturatingCounter_93_io_enable),
    .io_value(SaturatingCounter_93_io_value)
  );
  SaturatingCounter SaturatingCounter_94 (
    .clock(SaturatingCounter_94_clock),
    .reset(SaturatingCounter_94_reset),
    .io_enable(SaturatingCounter_94_io_enable),
    .io_value(SaturatingCounter_94_io_value)
  );
  SaturatingCounter SaturatingCounter_95 (
    .clock(SaturatingCounter_95_clock),
    .reset(SaturatingCounter_95_reset),
    .io_enable(SaturatingCounter_95_io_enable),
    .io_value(SaturatingCounter_95_io_value)
  );
  SaturatingCounter SaturatingCounter_96 (
    .clock(SaturatingCounter_96_clock),
    .reset(SaturatingCounter_96_reset),
    .io_enable(SaturatingCounter_96_io_enable),
    .io_value(SaturatingCounter_96_io_value)
  );
  SaturatingCounter SaturatingCounter_97 (
    .clock(SaturatingCounter_97_clock),
    .reset(SaturatingCounter_97_reset),
    .io_enable(SaturatingCounter_97_io_enable),
    .io_value(SaturatingCounter_97_io_value)
  );
  SaturatingCounter SaturatingCounter_98 (
    .clock(SaturatingCounter_98_clock),
    .reset(SaturatingCounter_98_reset),
    .io_enable(SaturatingCounter_98_io_enable),
    .io_value(SaturatingCounter_98_io_value)
  );
  SaturatingCounter SaturatingCounter_99 (
    .clock(SaturatingCounter_99_clock),
    .reset(SaturatingCounter_99_reset),
    .io_enable(SaturatingCounter_99_io_enable),
    .io_value(SaturatingCounter_99_io_value)
  );
  SaturatingCounter SaturatingCounter_100 (
    .clock(SaturatingCounter_100_clock),
    .reset(SaturatingCounter_100_reset),
    .io_enable(SaturatingCounter_100_io_enable),
    .io_value(SaturatingCounter_100_io_value)
  );
  SaturatingCounter SaturatingCounter_101 (
    .clock(SaturatingCounter_101_clock),
    .reset(SaturatingCounter_101_reset),
    .io_enable(SaturatingCounter_101_io_enable),
    .io_value(SaturatingCounter_101_io_value)
  );
  SaturatingCounter SaturatingCounter_102 (
    .clock(SaturatingCounter_102_clock),
    .reset(SaturatingCounter_102_reset),
    .io_enable(SaturatingCounter_102_io_enable),
    .io_value(SaturatingCounter_102_io_value)
  );
  SaturatingCounter SaturatingCounter_103 (
    .clock(SaturatingCounter_103_clock),
    .reset(SaturatingCounter_103_reset),
    .io_enable(SaturatingCounter_103_io_enable),
    .io_value(SaturatingCounter_103_io_value)
  );
  SaturatingCounter SaturatingCounter_104 (
    .clock(SaturatingCounter_104_clock),
    .reset(SaturatingCounter_104_reset),
    .io_enable(SaturatingCounter_104_io_enable),
    .io_value(SaturatingCounter_104_io_value)
  );
  SaturatingCounter SaturatingCounter_105 (
    .clock(SaturatingCounter_105_clock),
    .reset(SaturatingCounter_105_reset),
    .io_enable(SaturatingCounter_105_io_enable),
    .io_value(SaturatingCounter_105_io_value)
  );
  SaturatingCounter SaturatingCounter_106 (
    .clock(SaturatingCounter_106_clock),
    .reset(SaturatingCounter_106_reset),
    .io_enable(SaturatingCounter_106_io_enable),
    .io_value(SaturatingCounter_106_io_value)
  );
  SaturatingCounter SaturatingCounter_107 (
    .clock(SaturatingCounter_107_clock),
    .reset(SaturatingCounter_107_reset),
    .io_enable(SaturatingCounter_107_io_enable),
    .io_value(SaturatingCounter_107_io_value)
  );
  SaturatingCounter SaturatingCounter_108 (
    .clock(SaturatingCounter_108_clock),
    .reset(SaturatingCounter_108_reset),
    .io_enable(SaturatingCounter_108_io_enable),
    .io_value(SaturatingCounter_108_io_value)
  );
  SaturatingCounter SaturatingCounter_109 (
    .clock(SaturatingCounter_109_clock),
    .reset(SaturatingCounter_109_reset),
    .io_enable(SaturatingCounter_109_io_enable),
    .io_value(SaturatingCounter_109_io_value)
  );
  SaturatingCounter SaturatingCounter_110 (
    .clock(SaturatingCounter_110_clock),
    .reset(SaturatingCounter_110_reset),
    .io_enable(SaturatingCounter_110_io_enable),
    .io_value(SaturatingCounter_110_io_value)
  );
  SaturatingCounter SaturatingCounter_111 (
    .clock(SaturatingCounter_111_clock),
    .reset(SaturatingCounter_111_reset),
    .io_enable(SaturatingCounter_111_io_enable),
    .io_value(SaturatingCounter_111_io_value)
  );
  SaturatingCounter SaturatingCounter_112 (
    .clock(SaturatingCounter_112_clock),
    .reset(SaturatingCounter_112_reset),
    .io_enable(SaturatingCounter_112_io_enable),
    .io_value(SaturatingCounter_112_io_value)
  );
  SaturatingCounter SaturatingCounter_113 (
    .clock(SaturatingCounter_113_clock),
    .reset(SaturatingCounter_113_reset),
    .io_enable(SaturatingCounter_113_io_enable),
    .io_value(SaturatingCounter_113_io_value)
  );
  SaturatingCounter SaturatingCounter_114 (
    .clock(SaturatingCounter_114_clock),
    .reset(SaturatingCounter_114_reset),
    .io_enable(SaturatingCounter_114_io_enable),
    .io_value(SaturatingCounter_114_io_value)
  );
  SaturatingCounter SaturatingCounter_115 (
    .clock(SaturatingCounter_115_clock),
    .reset(SaturatingCounter_115_reset),
    .io_enable(SaturatingCounter_115_io_enable),
    .io_value(SaturatingCounter_115_io_value)
  );
  SaturatingCounter SaturatingCounter_116 (
    .clock(SaturatingCounter_116_clock),
    .reset(SaturatingCounter_116_reset),
    .io_enable(SaturatingCounter_116_io_enable),
    .io_value(SaturatingCounter_116_io_value)
  );
  SaturatingCounter SaturatingCounter_117 (
    .clock(SaturatingCounter_117_clock),
    .reset(SaturatingCounter_117_reset),
    .io_enable(SaturatingCounter_117_io_enable),
    .io_value(SaturatingCounter_117_io_value)
  );
  SaturatingCounter SaturatingCounter_118 (
    .clock(SaturatingCounter_118_clock),
    .reset(SaturatingCounter_118_reset),
    .io_enable(SaturatingCounter_118_io_enable),
    .io_value(SaturatingCounter_118_io_value)
  );
  SaturatingCounter SaturatingCounter_119 (
    .clock(SaturatingCounter_119_clock),
    .reset(SaturatingCounter_119_reset),
    .io_enable(SaturatingCounter_119_io_enable),
    .io_value(SaturatingCounter_119_io_value)
  );
  SaturatingCounter SaturatingCounter_120 (
    .clock(SaturatingCounter_120_clock),
    .reset(SaturatingCounter_120_reset),
    .io_enable(SaturatingCounter_120_io_enable),
    .io_value(SaturatingCounter_120_io_value)
  );
  SaturatingCounter SaturatingCounter_121 (
    .clock(SaturatingCounter_121_clock),
    .reset(SaturatingCounter_121_reset),
    .io_enable(SaturatingCounter_121_io_enable),
    .io_value(SaturatingCounter_121_io_value)
  );
  SaturatingCounter SaturatingCounter_122 (
    .clock(SaturatingCounter_122_clock),
    .reset(SaturatingCounter_122_reset),
    .io_enable(SaturatingCounter_122_io_enable),
    .io_value(SaturatingCounter_122_io_value)
  );
  SaturatingCounter SaturatingCounter_123 (
    .clock(SaturatingCounter_123_clock),
    .reset(SaturatingCounter_123_reset),
    .io_enable(SaturatingCounter_123_io_enable),
    .io_value(SaturatingCounter_123_io_value)
  );
  SaturatingCounter SaturatingCounter_124 (
    .clock(SaturatingCounter_124_clock),
    .reset(SaturatingCounter_124_reset),
    .io_enable(SaturatingCounter_124_io_enable),
    .io_value(SaturatingCounter_124_io_value)
  );
  SaturatingCounter SaturatingCounter_125 (
    .clock(SaturatingCounter_125_clock),
    .reset(SaturatingCounter_125_reset),
    .io_enable(SaturatingCounter_125_io_enable),
    .io_value(SaturatingCounter_125_io_value)
  );
  SaturatingCounter SaturatingCounter_126 (
    .clock(SaturatingCounter_126_clock),
    .reset(SaturatingCounter_126_reset),
    .io_enable(SaturatingCounter_126_io_enable),
    .io_value(SaturatingCounter_126_io_value)
  );
  SaturatingCounter SaturatingCounter_127 (
    .clock(SaturatingCounter_127_clock),
    .reset(SaturatingCounter_127_reset),
    .io_enable(SaturatingCounter_127_io_enable),
    .io_value(SaturatingCounter_127_io_value)
  );
  SaturatingCounter SaturatingCounter_128 (
    .clock(SaturatingCounter_128_clock),
    .reset(SaturatingCounter_128_reset),
    .io_enable(SaturatingCounter_128_io_enable),
    .io_value(SaturatingCounter_128_io_value)
  );
  SaturatingCounter SaturatingCounter_129 (
    .clock(SaturatingCounter_129_clock),
    .reset(SaturatingCounter_129_reset),
    .io_enable(SaturatingCounter_129_io_enable),
    .io_value(SaturatingCounter_129_io_value)
  );
  SaturatingCounter SaturatingCounter_130 (
    .clock(SaturatingCounter_130_clock),
    .reset(SaturatingCounter_130_reset),
    .io_enable(SaturatingCounter_130_io_enable),
    .io_value(SaturatingCounter_130_io_value)
  );
  SaturatingCounter SaturatingCounter_131 (
    .clock(SaturatingCounter_131_clock),
    .reset(SaturatingCounter_131_reset),
    .io_enable(SaturatingCounter_131_io_enable),
    .io_value(SaturatingCounter_131_io_value)
  );
  SaturatingCounter SaturatingCounter_132 (
    .clock(SaturatingCounter_132_clock),
    .reset(SaturatingCounter_132_reset),
    .io_enable(SaturatingCounter_132_io_enable),
    .io_value(SaturatingCounter_132_io_value)
  );
  SaturatingCounter SaturatingCounter_133 (
    .clock(SaturatingCounter_133_clock),
    .reset(SaturatingCounter_133_reset),
    .io_enable(SaturatingCounter_133_io_enable),
    .io_value(SaturatingCounter_133_io_value)
  );
  SaturatingCounter SaturatingCounter_134 (
    .clock(SaturatingCounter_134_clock),
    .reset(SaturatingCounter_134_reset),
    .io_enable(SaturatingCounter_134_io_enable),
    .io_value(SaturatingCounter_134_io_value)
  );
  SaturatingCounter SaturatingCounter_135 (
    .clock(SaturatingCounter_135_clock),
    .reset(SaturatingCounter_135_reset),
    .io_enable(SaturatingCounter_135_io_enable),
    .io_value(SaturatingCounter_135_io_value)
  );
  SaturatingCounter SaturatingCounter_136 (
    .clock(SaturatingCounter_136_clock),
    .reset(SaturatingCounter_136_reset),
    .io_enable(SaturatingCounter_136_io_enable),
    .io_value(SaturatingCounter_136_io_value)
  );
  SaturatingCounter SaturatingCounter_137 (
    .clock(SaturatingCounter_137_clock),
    .reset(SaturatingCounter_137_reset),
    .io_enable(SaturatingCounter_137_io_enable),
    .io_value(SaturatingCounter_137_io_value)
  );
  SaturatingCounter SaturatingCounter_138 (
    .clock(SaturatingCounter_138_clock),
    .reset(SaturatingCounter_138_reset),
    .io_enable(SaturatingCounter_138_io_enable),
    .io_value(SaturatingCounter_138_io_value)
  );
  SaturatingCounter SaturatingCounter_139 (
    .clock(SaturatingCounter_139_clock),
    .reset(SaturatingCounter_139_reset),
    .io_enable(SaturatingCounter_139_io_enable),
    .io_value(SaturatingCounter_139_io_value)
  );
  SaturatingCounter SaturatingCounter_140 (
    .clock(SaturatingCounter_140_clock),
    .reset(SaturatingCounter_140_reset),
    .io_enable(SaturatingCounter_140_io_enable),
    .io_value(SaturatingCounter_140_io_value)
  );
  SaturatingCounter SaturatingCounter_141 (
    .clock(SaturatingCounter_141_clock),
    .reset(SaturatingCounter_141_reset),
    .io_enable(SaturatingCounter_141_io_enable),
    .io_value(SaturatingCounter_141_io_value)
  );
  SaturatingCounter SaturatingCounter_142 (
    .clock(SaturatingCounter_142_clock),
    .reset(SaturatingCounter_142_reset),
    .io_enable(SaturatingCounter_142_io_enable),
    .io_value(SaturatingCounter_142_io_value)
  );
  SaturatingCounter SaturatingCounter_143 (
    .clock(SaturatingCounter_143_clock),
    .reset(SaturatingCounter_143_reset),
    .io_enable(SaturatingCounter_143_io_enable),
    .io_value(SaturatingCounter_143_io_value)
  );
  SaturatingCounter SaturatingCounter_144 (
    .clock(SaturatingCounter_144_clock),
    .reset(SaturatingCounter_144_reset),
    .io_enable(SaturatingCounter_144_io_enable),
    .io_value(SaturatingCounter_144_io_value)
  );
  SaturatingCounter SaturatingCounter_145 (
    .clock(SaturatingCounter_145_clock),
    .reset(SaturatingCounter_145_reset),
    .io_enable(SaturatingCounter_145_io_enable),
    .io_value(SaturatingCounter_145_io_value)
  );
  SaturatingCounter SaturatingCounter_146 (
    .clock(SaturatingCounter_146_clock),
    .reset(SaturatingCounter_146_reset),
    .io_enable(SaturatingCounter_146_io_enable),
    .io_value(SaturatingCounter_146_io_value)
  );
  SaturatingCounter SaturatingCounter_147 (
    .clock(SaturatingCounter_147_clock),
    .reset(SaturatingCounter_147_reset),
    .io_enable(SaturatingCounter_147_io_enable),
    .io_value(SaturatingCounter_147_io_value)
  );
  SaturatingCounter SaturatingCounter_148 (
    .clock(SaturatingCounter_148_clock),
    .reset(SaturatingCounter_148_reset),
    .io_enable(SaturatingCounter_148_io_enable),
    .io_value(SaturatingCounter_148_io_value)
  );
  SaturatingCounter SaturatingCounter_149 (
    .clock(SaturatingCounter_149_clock),
    .reset(SaturatingCounter_149_reset),
    .io_enable(SaturatingCounter_149_io_enable),
    .io_value(SaturatingCounter_149_io_value)
  );
  SaturatingCounter SaturatingCounter_150 (
    .clock(SaturatingCounter_150_clock),
    .reset(SaturatingCounter_150_reset),
    .io_enable(SaturatingCounter_150_io_enable),
    .io_value(SaturatingCounter_150_io_value)
  );
  SaturatingCounter SaturatingCounter_151 (
    .clock(SaturatingCounter_151_clock),
    .reset(SaturatingCounter_151_reset),
    .io_enable(SaturatingCounter_151_io_enable),
    .io_value(SaturatingCounter_151_io_value)
  );
  SaturatingCounter SaturatingCounter_152 (
    .clock(SaturatingCounter_152_clock),
    .reset(SaturatingCounter_152_reset),
    .io_enable(SaturatingCounter_152_io_enable),
    .io_value(SaturatingCounter_152_io_value)
  );
  SaturatingCounter SaturatingCounter_153 (
    .clock(SaturatingCounter_153_clock),
    .reset(SaturatingCounter_153_reset),
    .io_enable(SaturatingCounter_153_io_enable),
    .io_value(SaturatingCounter_153_io_value)
  );
  SaturatingCounter SaturatingCounter_154 (
    .clock(SaturatingCounter_154_clock),
    .reset(SaturatingCounter_154_reset),
    .io_enable(SaturatingCounter_154_io_enable),
    .io_value(SaturatingCounter_154_io_value)
  );
  SaturatingCounter SaturatingCounter_155 (
    .clock(SaturatingCounter_155_clock),
    .reset(SaturatingCounter_155_reset),
    .io_enable(SaturatingCounter_155_io_enable),
    .io_value(SaturatingCounter_155_io_value)
  );
  SaturatingCounter SaturatingCounter_156 (
    .clock(SaturatingCounter_156_clock),
    .reset(SaturatingCounter_156_reset),
    .io_enable(SaturatingCounter_156_io_enable),
    .io_value(SaturatingCounter_156_io_value)
  );
  SaturatingCounter SaturatingCounter_157 (
    .clock(SaturatingCounter_157_clock),
    .reset(SaturatingCounter_157_reset),
    .io_enable(SaturatingCounter_157_io_enable),
    .io_value(SaturatingCounter_157_io_value)
  );
  SaturatingCounter SaturatingCounter_158 (
    .clock(SaturatingCounter_158_clock),
    .reset(SaturatingCounter_158_reset),
    .io_enable(SaturatingCounter_158_io_enable),
    .io_value(SaturatingCounter_158_io_value)
  );
  SaturatingCounter SaturatingCounter_159 (
    .clock(SaturatingCounter_159_clock),
    .reset(SaturatingCounter_159_reset),
    .io_enable(SaturatingCounter_159_io_enable),
    .io_value(SaturatingCounter_159_io_value)
  );
  SaturatingCounter SaturatingCounter_160 (
    .clock(SaturatingCounter_160_clock),
    .reset(SaturatingCounter_160_reset),
    .io_enable(SaturatingCounter_160_io_enable),
    .io_value(SaturatingCounter_160_io_value)
  );
  SaturatingCounter SaturatingCounter_161 (
    .clock(SaturatingCounter_161_clock),
    .reset(SaturatingCounter_161_reset),
    .io_enable(SaturatingCounter_161_io_enable),
    .io_value(SaturatingCounter_161_io_value)
  );
  SaturatingCounter SaturatingCounter_162 (
    .clock(SaturatingCounter_162_clock),
    .reset(SaturatingCounter_162_reset),
    .io_enable(SaturatingCounter_162_io_enable),
    .io_value(SaturatingCounter_162_io_value)
  );
  SaturatingCounter SaturatingCounter_163 (
    .clock(SaturatingCounter_163_clock),
    .reset(SaturatingCounter_163_reset),
    .io_enable(SaturatingCounter_163_io_enable),
    .io_value(SaturatingCounter_163_io_value)
  );
  SaturatingCounter SaturatingCounter_164 (
    .clock(SaturatingCounter_164_clock),
    .reset(SaturatingCounter_164_reset),
    .io_enable(SaturatingCounter_164_io_enable),
    .io_value(SaturatingCounter_164_io_value)
  );
  SaturatingCounter SaturatingCounter_165 (
    .clock(SaturatingCounter_165_clock),
    .reset(SaturatingCounter_165_reset),
    .io_enable(SaturatingCounter_165_io_enable),
    .io_value(SaturatingCounter_165_io_value)
  );
  SaturatingCounter SaturatingCounter_166 (
    .clock(SaturatingCounter_166_clock),
    .reset(SaturatingCounter_166_reset),
    .io_enable(SaturatingCounter_166_io_enable),
    .io_value(SaturatingCounter_166_io_value)
  );
  SaturatingCounter SaturatingCounter_167 (
    .clock(SaturatingCounter_167_clock),
    .reset(SaturatingCounter_167_reset),
    .io_enable(SaturatingCounter_167_io_enable),
    .io_value(SaturatingCounter_167_io_value)
  );
  SaturatingCounter SaturatingCounter_168 (
    .clock(SaturatingCounter_168_clock),
    .reset(SaturatingCounter_168_reset),
    .io_enable(SaturatingCounter_168_io_enable),
    .io_value(SaturatingCounter_168_io_value)
  );
  SaturatingCounter SaturatingCounter_169 (
    .clock(SaturatingCounter_169_clock),
    .reset(SaturatingCounter_169_reset),
    .io_enable(SaturatingCounter_169_io_enable),
    .io_value(SaturatingCounter_169_io_value)
  );
  SaturatingCounter SaturatingCounter_170 (
    .clock(SaturatingCounter_170_clock),
    .reset(SaturatingCounter_170_reset),
    .io_enable(SaturatingCounter_170_io_enable),
    .io_value(SaturatingCounter_170_io_value)
  );
  SaturatingCounter SaturatingCounter_171 (
    .clock(SaturatingCounter_171_clock),
    .reset(SaturatingCounter_171_reset),
    .io_enable(SaturatingCounter_171_io_enable),
    .io_value(SaturatingCounter_171_io_value)
  );
  SaturatingCounter SaturatingCounter_172 (
    .clock(SaturatingCounter_172_clock),
    .reset(SaturatingCounter_172_reset),
    .io_enable(SaturatingCounter_172_io_enable),
    .io_value(SaturatingCounter_172_io_value)
  );
  SaturatingCounter SaturatingCounter_173 (
    .clock(SaturatingCounter_173_clock),
    .reset(SaturatingCounter_173_reset),
    .io_enable(SaturatingCounter_173_io_enable),
    .io_value(SaturatingCounter_173_io_value)
  );
  SaturatingCounter SaturatingCounter_174 (
    .clock(SaturatingCounter_174_clock),
    .reset(SaturatingCounter_174_reset),
    .io_enable(SaturatingCounter_174_io_enable),
    .io_value(SaturatingCounter_174_io_value)
  );
  SaturatingCounter SaturatingCounter_175 (
    .clock(SaturatingCounter_175_clock),
    .reset(SaturatingCounter_175_reset),
    .io_enable(SaturatingCounter_175_io_enable),
    .io_value(SaturatingCounter_175_io_value)
  );
  SaturatingCounter SaturatingCounter_176 (
    .clock(SaturatingCounter_176_clock),
    .reset(SaturatingCounter_176_reset),
    .io_enable(SaturatingCounter_176_io_enable),
    .io_value(SaturatingCounter_176_io_value)
  );
  SaturatingCounter SaturatingCounter_177 (
    .clock(SaturatingCounter_177_clock),
    .reset(SaturatingCounter_177_reset),
    .io_enable(SaturatingCounter_177_io_enable),
    .io_value(SaturatingCounter_177_io_value)
  );
  SaturatingCounter SaturatingCounter_178 (
    .clock(SaturatingCounter_178_clock),
    .reset(SaturatingCounter_178_reset),
    .io_enable(SaturatingCounter_178_io_enable),
    .io_value(SaturatingCounter_178_io_value)
  );
  SaturatingCounter SaturatingCounter_179 (
    .clock(SaturatingCounter_179_clock),
    .reset(SaturatingCounter_179_reset),
    .io_enable(SaturatingCounter_179_io_enable),
    .io_value(SaturatingCounter_179_io_value)
  );
  SaturatingCounter SaturatingCounter_180 (
    .clock(SaturatingCounter_180_clock),
    .reset(SaturatingCounter_180_reset),
    .io_enable(SaturatingCounter_180_io_enable),
    .io_value(SaturatingCounter_180_io_value)
  );
  SaturatingCounter SaturatingCounter_181 (
    .clock(SaturatingCounter_181_clock),
    .reset(SaturatingCounter_181_reset),
    .io_enable(SaturatingCounter_181_io_enable),
    .io_value(SaturatingCounter_181_io_value)
  );
  SaturatingCounter SaturatingCounter_182 (
    .clock(SaturatingCounter_182_clock),
    .reset(SaturatingCounter_182_reset),
    .io_enable(SaturatingCounter_182_io_enable),
    .io_value(SaturatingCounter_182_io_value)
  );
  SaturatingCounter SaturatingCounter_183 (
    .clock(SaturatingCounter_183_clock),
    .reset(SaturatingCounter_183_reset),
    .io_enable(SaturatingCounter_183_io_enable),
    .io_value(SaturatingCounter_183_io_value)
  );
  SaturatingCounter SaturatingCounter_184 (
    .clock(SaturatingCounter_184_clock),
    .reset(SaturatingCounter_184_reset),
    .io_enable(SaturatingCounter_184_io_enable),
    .io_value(SaturatingCounter_184_io_value)
  );
  SaturatingCounter SaturatingCounter_185 (
    .clock(SaturatingCounter_185_clock),
    .reset(SaturatingCounter_185_reset),
    .io_enable(SaturatingCounter_185_io_enable),
    .io_value(SaturatingCounter_185_io_value)
  );
  SaturatingCounter SaturatingCounter_186 (
    .clock(SaturatingCounter_186_clock),
    .reset(SaturatingCounter_186_reset),
    .io_enable(SaturatingCounter_186_io_enable),
    .io_value(SaturatingCounter_186_io_value)
  );
  SaturatingCounter SaturatingCounter_187 (
    .clock(SaturatingCounter_187_clock),
    .reset(SaturatingCounter_187_reset),
    .io_enable(SaturatingCounter_187_io_enable),
    .io_value(SaturatingCounter_187_io_value)
  );
  SaturatingCounter SaturatingCounter_188 (
    .clock(SaturatingCounter_188_clock),
    .reset(SaturatingCounter_188_reset),
    .io_enable(SaturatingCounter_188_io_enable),
    .io_value(SaturatingCounter_188_io_value)
  );
  SaturatingCounter SaturatingCounter_189 (
    .clock(SaturatingCounter_189_clock),
    .reset(SaturatingCounter_189_reset),
    .io_enable(SaturatingCounter_189_io_enable),
    .io_value(SaturatingCounter_189_io_value)
  );
  SaturatingCounter SaturatingCounter_190 (
    .clock(SaturatingCounter_190_clock),
    .reset(SaturatingCounter_190_reset),
    .io_enable(SaturatingCounter_190_io_enable),
    .io_value(SaturatingCounter_190_io_value)
  );
  SaturatingCounter SaturatingCounter_191 (
    .clock(SaturatingCounter_191_clock),
    .reset(SaturatingCounter_191_reset),
    .io_enable(SaturatingCounter_191_io_enable),
    .io_value(SaturatingCounter_191_io_value)
  );
  SaturatingCounter SaturatingCounter_192 (
    .clock(SaturatingCounter_192_clock),
    .reset(SaturatingCounter_192_reset),
    .io_enable(SaturatingCounter_192_io_enable),
    .io_value(SaturatingCounter_192_io_value)
  );
  SaturatingCounter SaturatingCounter_193 (
    .clock(SaturatingCounter_193_clock),
    .reset(SaturatingCounter_193_reset),
    .io_enable(SaturatingCounter_193_io_enable),
    .io_value(SaturatingCounter_193_io_value)
  );
  SaturatingCounter SaturatingCounter_194 (
    .clock(SaturatingCounter_194_clock),
    .reset(SaturatingCounter_194_reset),
    .io_enable(SaturatingCounter_194_io_enable),
    .io_value(SaturatingCounter_194_io_value)
  );
  SaturatingCounter SaturatingCounter_195 (
    .clock(SaturatingCounter_195_clock),
    .reset(SaturatingCounter_195_reset),
    .io_enable(SaturatingCounter_195_io_enable),
    .io_value(SaturatingCounter_195_io_value)
  );
  SaturatingCounter SaturatingCounter_196 (
    .clock(SaturatingCounter_196_clock),
    .reset(SaturatingCounter_196_reset),
    .io_enable(SaturatingCounter_196_io_enable),
    .io_value(SaturatingCounter_196_io_value)
  );
  SaturatingCounter SaturatingCounter_197 (
    .clock(SaturatingCounter_197_clock),
    .reset(SaturatingCounter_197_reset),
    .io_enable(SaturatingCounter_197_io_enable),
    .io_value(SaturatingCounter_197_io_value)
  );
  SaturatingCounter SaturatingCounter_198 (
    .clock(SaturatingCounter_198_clock),
    .reset(SaturatingCounter_198_reset),
    .io_enable(SaturatingCounter_198_io_enable),
    .io_value(SaturatingCounter_198_io_value)
  );
  SaturatingCounter SaturatingCounter_199 (
    .clock(SaturatingCounter_199_clock),
    .reset(SaturatingCounter_199_reset),
    .io_enable(SaturatingCounter_199_io_enable),
    .io_value(SaturatingCounter_199_io_value)
  );
  SaturatingCounter SaturatingCounter_200 (
    .clock(SaturatingCounter_200_clock),
    .reset(SaturatingCounter_200_reset),
    .io_enable(SaturatingCounter_200_io_enable),
    .io_value(SaturatingCounter_200_io_value)
  );
  SaturatingCounter SaturatingCounter_201 (
    .clock(SaturatingCounter_201_clock),
    .reset(SaturatingCounter_201_reset),
    .io_enable(SaturatingCounter_201_io_enable),
    .io_value(SaturatingCounter_201_io_value)
  );
  SaturatingCounter SaturatingCounter_202 (
    .clock(SaturatingCounter_202_clock),
    .reset(SaturatingCounter_202_reset),
    .io_enable(SaturatingCounter_202_io_enable),
    .io_value(SaturatingCounter_202_io_value)
  );
  SaturatingCounter SaturatingCounter_203 (
    .clock(SaturatingCounter_203_clock),
    .reset(SaturatingCounter_203_reset),
    .io_enable(SaturatingCounter_203_io_enable),
    .io_value(SaturatingCounter_203_io_value)
  );
  SaturatingCounter SaturatingCounter_204 (
    .clock(SaturatingCounter_204_clock),
    .reset(SaturatingCounter_204_reset),
    .io_enable(SaturatingCounter_204_io_enable),
    .io_value(SaturatingCounter_204_io_value)
  );
  SaturatingCounter SaturatingCounter_205 (
    .clock(SaturatingCounter_205_clock),
    .reset(SaturatingCounter_205_reset),
    .io_enable(SaturatingCounter_205_io_enable),
    .io_value(SaturatingCounter_205_io_value)
  );
  SaturatingCounter SaturatingCounter_206 (
    .clock(SaturatingCounter_206_clock),
    .reset(SaturatingCounter_206_reset),
    .io_enable(SaturatingCounter_206_io_enable),
    .io_value(SaturatingCounter_206_io_value)
  );
  SaturatingCounter SaturatingCounter_207 (
    .clock(SaturatingCounter_207_clock),
    .reset(SaturatingCounter_207_reset),
    .io_enable(SaturatingCounter_207_io_enable),
    .io_value(SaturatingCounter_207_io_value)
  );
  SaturatingCounter SaturatingCounter_208 (
    .clock(SaturatingCounter_208_clock),
    .reset(SaturatingCounter_208_reset),
    .io_enable(SaturatingCounter_208_io_enable),
    .io_value(SaturatingCounter_208_io_value)
  );
  SaturatingCounter SaturatingCounter_209 (
    .clock(SaturatingCounter_209_clock),
    .reset(SaturatingCounter_209_reset),
    .io_enable(SaturatingCounter_209_io_enable),
    .io_value(SaturatingCounter_209_io_value)
  );
  SaturatingCounter SaturatingCounter_210 (
    .clock(SaturatingCounter_210_clock),
    .reset(SaturatingCounter_210_reset),
    .io_enable(SaturatingCounter_210_io_enable),
    .io_value(SaturatingCounter_210_io_value)
  );
  SaturatingCounter SaturatingCounter_211 (
    .clock(SaturatingCounter_211_clock),
    .reset(SaturatingCounter_211_reset),
    .io_enable(SaturatingCounter_211_io_enable),
    .io_value(SaturatingCounter_211_io_value)
  );
  SaturatingCounter SaturatingCounter_212 (
    .clock(SaturatingCounter_212_clock),
    .reset(SaturatingCounter_212_reset),
    .io_enable(SaturatingCounter_212_io_enable),
    .io_value(SaturatingCounter_212_io_value)
  );
  SaturatingCounter SaturatingCounter_213 (
    .clock(SaturatingCounter_213_clock),
    .reset(SaturatingCounter_213_reset),
    .io_enable(SaturatingCounter_213_io_enable),
    .io_value(SaturatingCounter_213_io_value)
  );
  SaturatingCounter SaturatingCounter_214 (
    .clock(SaturatingCounter_214_clock),
    .reset(SaturatingCounter_214_reset),
    .io_enable(SaturatingCounter_214_io_enable),
    .io_value(SaturatingCounter_214_io_value)
  );
  SaturatingCounter SaturatingCounter_215 (
    .clock(SaturatingCounter_215_clock),
    .reset(SaturatingCounter_215_reset),
    .io_enable(SaturatingCounter_215_io_enable),
    .io_value(SaturatingCounter_215_io_value)
  );
  SaturatingCounter SaturatingCounter_216 (
    .clock(SaturatingCounter_216_clock),
    .reset(SaturatingCounter_216_reset),
    .io_enable(SaturatingCounter_216_io_enable),
    .io_value(SaturatingCounter_216_io_value)
  );
  SaturatingCounter SaturatingCounter_217 (
    .clock(SaturatingCounter_217_clock),
    .reset(SaturatingCounter_217_reset),
    .io_enable(SaturatingCounter_217_io_enable),
    .io_value(SaturatingCounter_217_io_value)
  );
  SaturatingCounter SaturatingCounter_218 (
    .clock(SaturatingCounter_218_clock),
    .reset(SaturatingCounter_218_reset),
    .io_enable(SaturatingCounter_218_io_enable),
    .io_value(SaturatingCounter_218_io_value)
  );
  SaturatingCounter SaturatingCounter_219 (
    .clock(SaturatingCounter_219_clock),
    .reset(SaturatingCounter_219_reset),
    .io_enable(SaturatingCounter_219_io_enable),
    .io_value(SaturatingCounter_219_io_value)
  );
  SaturatingCounter SaturatingCounter_220 (
    .clock(SaturatingCounter_220_clock),
    .reset(SaturatingCounter_220_reset),
    .io_enable(SaturatingCounter_220_io_enable),
    .io_value(SaturatingCounter_220_io_value)
  );
  SaturatingCounter SaturatingCounter_221 (
    .clock(SaturatingCounter_221_clock),
    .reset(SaturatingCounter_221_reset),
    .io_enable(SaturatingCounter_221_io_enable),
    .io_value(SaturatingCounter_221_io_value)
  );
  SaturatingCounter SaturatingCounter_222 (
    .clock(SaturatingCounter_222_clock),
    .reset(SaturatingCounter_222_reset),
    .io_enable(SaturatingCounter_222_io_enable),
    .io_value(SaturatingCounter_222_io_value)
  );
  SaturatingCounter SaturatingCounter_223 (
    .clock(SaturatingCounter_223_clock),
    .reset(SaturatingCounter_223_reset),
    .io_enable(SaturatingCounter_223_io_enable),
    .io_value(SaturatingCounter_223_io_value)
  );
  SaturatingCounter SaturatingCounter_224 (
    .clock(SaturatingCounter_224_clock),
    .reset(SaturatingCounter_224_reset),
    .io_enable(SaturatingCounter_224_io_enable),
    .io_value(SaturatingCounter_224_io_value)
  );
  SaturatingCounter SaturatingCounter_225 (
    .clock(SaturatingCounter_225_clock),
    .reset(SaturatingCounter_225_reset),
    .io_enable(SaturatingCounter_225_io_enable),
    .io_value(SaturatingCounter_225_io_value)
  );
  SaturatingCounter SaturatingCounter_226 (
    .clock(SaturatingCounter_226_clock),
    .reset(SaturatingCounter_226_reset),
    .io_enable(SaturatingCounter_226_io_enable),
    .io_value(SaturatingCounter_226_io_value)
  );
  SaturatingCounter SaturatingCounter_227 (
    .clock(SaturatingCounter_227_clock),
    .reset(SaturatingCounter_227_reset),
    .io_enable(SaturatingCounter_227_io_enable),
    .io_value(SaturatingCounter_227_io_value)
  );
  SaturatingCounter SaturatingCounter_228 (
    .clock(SaturatingCounter_228_clock),
    .reset(SaturatingCounter_228_reset),
    .io_enable(SaturatingCounter_228_io_enable),
    .io_value(SaturatingCounter_228_io_value)
  );
  SaturatingCounter SaturatingCounter_229 (
    .clock(SaturatingCounter_229_clock),
    .reset(SaturatingCounter_229_reset),
    .io_enable(SaturatingCounter_229_io_enable),
    .io_value(SaturatingCounter_229_io_value)
  );
  SaturatingCounter SaturatingCounter_230 (
    .clock(SaturatingCounter_230_clock),
    .reset(SaturatingCounter_230_reset),
    .io_enable(SaturatingCounter_230_io_enable),
    .io_value(SaturatingCounter_230_io_value)
  );
  SaturatingCounter SaturatingCounter_231 (
    .clock(SaturatingCounter_231_clock),
    .reset(SaturatingCounter_231_reset),
    .io_enable(SaturatingCounter_231_io_enable),
    .io_value(SaturatingCounter_231_io_value)
  );
  SaturatingCounter SaturatingCounter_232 (
    .clock(SaturatingCounter_232_clock),
    .reset(SaturatingCounter_232_reset),
    .io_enable(SaturatingCounter_232_io_enable),
    .io_value(SaturatingCounter_232_io_value)
  );
  SaturatingCounter SaturatingCounter_233 (
    .clock(SaturatingCounter_233_clock),
    .reset(SaturatingCounter_233_reset),
    .io_enable(SaturatingCounter_233_io_enable),
    .io_value(SaturatingCounter_233_io_value)
  );
  SaturatingCounter SaturatingCounter_234 (
    .clock(SaturatingCounter_234_clock),
    .reset(SaturatingCounter_234_reset),
    .io_enable(SaturatingCounter_234_io_enable),
    .io_value(SaturatingCounter_234_io_value)
  );
  SaturatingCounter SaturatingCounter_235 (
    .clock(SaturatingCounter_235_clock),
    .reset(SaturatingCounter_235_reset),
    .io_enable(SaturatingCounter_235_io_enable),
    .io_value(SaturatingCounter_235_io_value)
  );
  SaturatingCounter SaturatingCounter_236 (
    .clock(SaturatingCounter_236_clock),
    .reset(SaturatingCounter_236_reset),
    .io_enable(SaturatingCounter_236_io_enable),
    .io_value(SaturatingCounter_236_io_value)
  );
  SaturatingCounter SaturatingCounter_237 (
    .clock(SaturatingCounter_237_clock),
    .reset(SaturatingCounter_237_reset),
    .io_enable(SaturatingCounter_237_io_enable),
    .io_value(SaturatingCounter_237_io_value)
  );
  SaturatingCounter SaturatingCounter_238 (
    .clock(SaturatingCounter_238_clock),
    .reset(SaturatingCounter_238_reset),
    .io_enable(SaturatingCounter_238_io_enable),
    .io_value(SaturatingCounter_238_io_value)
  );
  SaturatingCounter SaturatingCounter_239 (
    .clock(SaturatingCounter_239_clock),
    .reset(SaturatingCounter_239_reset),
    .io_enable(SaturatingCounter_239_io_enable),
    .io_value(SaturatingCounter_239_io_value)
  );
  SaturatingCounter SaturatingCounter_240 (
    .clock(SaturatingCounter_240_clock),
    .reset(SaturatingCounter_240_reset),
    .io_enable(SaturatingCounter_240_io_enable),
    .io_value(SaturatingCounter_240_io_value)
  );
  SaturatingCounter SaturatingCounter_241 (
    .clock(SaturatingCounter_241_clock),
    .reset(SaturatingCounter_241_reset),
    .io_enable(SaturatingCounter_241_io_enable),
    .io_value(SaturatingCounter_241_io_value)
  );
  SaturatingCounter SaturatingCounter_242 (
    .clock(SaturatingCounter_242_clock),
    .reset(SaturatingCounter_242_reset),
    .io_enable(SaturatingCounter_242_io_enable),
    .io_value(SaturatingCounter_242_io_value)
  );
  SaturatingCounter SaturatingCounter_243 (
    .clock(SaturatingCounter_243_clock),
    .reset(SaturatingCounter_243_reset),
    .io_enable(SaturatingCounter_243_io_enable),
    .io_value(SaturatingCounter_243_io_value)
  );
  SaturatingCounter SaturatingCounter_244 (
    .clock(SaturatingCounter_244_clock),
    .reset(SaturatingCounter_244_reset),
    .io_enable(SaturatingCounter_244_io_enable),
    .io_value(SaturatingCounter_244_io_value)
  );
  SaturatingCounter SaturatingCounter_245 (
    .clock(SaturatingCounter_245_clock),
    .reset(SaturatingCounter_245_reset),
    .io_enable(SaturatingCounter_245_io_enable),
    .io_value(SaturatingCounter_245_io_value)
  );
  SaturatingCounter SaturatingCounter_246 (
    .clock(SaturatingCounter_246_clock),
    .reset(SaturatingCounter_246_reset),
    .io_enable(SaturatingCounter_246_io_enable),
    .io_value(SaturatingCounter_246_io_value)
  );
  SaturatingCounter SaturatingCounter_247 (
    .clock(SaturatingCounter_247_clock),
    .reset(SaturatingCounter_247_reset),
    .io_enable(SaturatingCounter_247_io_enable),
    .io_value(SaturatingCounter_247_io_value)
  );
  SaturatingCounter SaturatingCounter_248 (
    .clock(SaturatingCounter_248_clock),
    .reset(SaturatingCounter_248_reset),
    .io_enable(SaturatingCounter_248_io_enable),
    .io_value(SaturatingCounter_248_io_value)
  );
  SaturatingCounter SaturatingCounter_249 (
    .clock(SaturatingCounter_249_clock),
    .reset(SaturatingCounter_249_reset),
    .io_enable(SaturatingCounter_249_io_enable),
    .io_value(SaturatingCounter_249_io_value)
  );
  SaturatingCounter SaturatingCounter_250 (
    .clock(SaturatingCounter_250_clock),
    .reset(SaturatingCounter_250_reset),
    .io_enable(SaturatingCounter_250_io_enable),
    .io_value(SaturatingCounter_250_io_value)
  );
  SaturatingCounter SaturatingCounter_251 (
    .clock(SaturatingCounter_251_clock),
    .reset(SaturatingCounter_251_reset),
    .io_enable(SaturatingCounter_251_io_enable),
    .io_value(SaturatingCounter_251_io_value)
  );
  SaturatingCounter SaturatingCounter_252 (
    .clock(SaturatingCounter_252_clock),
    .reset(SaturatingCounter_252_reset),
    .io_enable(SaturatingCounter_252_io_enable),
    .io_value(SaturatingCounter_252_io_value)
  );
  SaturatingCounter SaturatingCounter_253 (
    .clock(SaturatingCounter_253_clock),
    .reset(SaturatingCounter_253_reset),
    .io_enable(SaturatingCounter_253_io_enable),
    .io_value(SaturatingCounter_253_io_value)
  );
  SaturatingCounter SaturatingCounter_254 (
    .clock(SaturatingCounter_254_clock),
    .reset(SaturatingCounter_254_reset),
    .io_enable(SaturatingCounter_254_io_enable),
    .io_value(SaturatingCounter_254_io_value)
  );
  SaturatingCounter SaturatingCounter_255 (
    .clock(SaturatingCounter_255_clock),
    .reset(SaturatingCounter_255_reset),
    .io_enable(SaturatingCounter_255_io_enable),
    .io_value(SaturatingCounter_255_io_value)
  );
  SaturatingCounter SaturatingCounter_256 (
    .clock(SaturatingCounter_256_clock),
    .reset(SaturatingCounter_256_reset),
    .io_enable(SaturatingCounter_256_io_enable),
    .io_value(SaturatingCounter_256_io_value)
  );
  SaturatingCounter SaturatingCounter_257 (
    .clock(SaturatingCounter_257_clock),
    .reset(SaturatingCounter_257_reset),
    .io_enable(SaturatingCounter_257_io_enable),
    .io_value(SaturatingCounter_257_io_value)
  );
  SaturatingCounter SaturatingCounter_258 (
    .clock(SaturatingCounter_258_clock),
    .reset(SaturatingCounter_258_reset),
    .io_enable(SaturatingCounter_258_io_enable),
    .io_value(SaturatingCounter_258_io_value)
  );
  SaturatingCounter SaturatingCounter_259 (
    .clock(SaturatingCounter_259_clock),
    .reset(SaturatingCounter_259_reset),
    .io_enable(SaturatingCounter_259_io_enable),
    .io_value(SaturatingCounter_259_io_value)
  );
  SaturatingCounter SaturatingCounter_260 (
    .clock(SaturatingCounter_260_clock),
    .reset(SaturatingCounter_260_reset),
    .io_enable(SaturatingCounter_260_io_enable),
    .io_value(SaturatingCounter_260_io_value)
  );
  SaturatingCounter SaturatingCounter_261 (
    .clock(SaturatingCounter_261_clock),
    .reset(SaturatingCounter_261_reset),
    .io_enable(SaturatingCounter_261_io_enable),
    .io_value(SaturatingCounter_261_io_value)
  );
  SaturatingCounter SaturatingCounter_262 (
    .clock(SaturatingCounter_262_clock),
    .reset(SaturatingCounter_262_reset),
    .io_enable(SaturatingCounter_262_io_enable),
    .io_value(SaturatingCounter_262_io_value)
  );
  SaturatingCounter SaturatingCounter_263 (
    .clock(SaturatingCounter_263_clock),
    .reset(SaturatingCounter_263_reset),
    .io_enable(SaturatingCounter_263_io_enable),
    .io_value(SaturatingCounter_263_io_value)
  );
  SaturatingCounter SaturatingCounter_264 (
    .clock(SaturatingCounter_264_clock),
    .reset(SaturatingCounter_264_reset),
    .io_enable(SaturatingCounter_264_io_enable),
    .io_value(SaturatingCounter_264_io_value)
  );
  SaturatingCounter SaturatingCounter_265 (
    .clock(SaturatingCounter_265_clock),
    .reset(SaturatingCounter_265_reset),
    .io_enable(SaturatingCounter_265_io_enable),
    .io_value(SaturatingCounter_265_io_value)
  );
  SaturatingCounter SaturatingCounter_266 (
    .clock(SaturatingCounter_266_clock),
    .reset(SaturatingCounter_266_reset),
    .io_enable(SaturatingCounter_266_io_enable),
    .io_value(SaturatingCounter_266_io_value)
  );
  SaturatingCounter SaturatingCounter_267 (
    .clock(SaturatingCounter_267_clock),
    .reset(SaturatingCounter_267_reset),
    .io_enable(SaturatingCounter_267_io_enable),
    .io_value(SaturatingCounter_267_io_value)
  );
  SaturatingCounter SaturatingCounter_268 (
    .clock(SaturatingCounter_268_clock),
    .reset(SaturatingCounter_268_reset),
    .io_enable(SaturatingCounter_268_io_enable),
    .io_value(SaturatingCounter_268_io_value)
  );
  SaturatingCounter SaturatingCounter_269 (
    .clock(SaturatingCounter_269_clock),
    .reset(SaturatingCounter_269_reset),
    .io_enable(SaturatingCounter_269_io_enable),
    .io_value(SaturatingCounter_269_io_value)
  );
  SaturatingCounter SaturatingCounter_270 (
    .clock(SaturatingCounter_270_clock),
    .reset(SaturatingCounter_270_reset),
    .io_enable(SaturatingCounter_270_io_enable),
    .io_value(SaturatingCounter_270_io_value)
  );
  SaturatingCounter SaturatingCounter_271 (
    .clock(SaturatingCounter_271_clock),
    .reset(SaturatingCounter_271_reset),
    .io_enable(SaturatingCounter_271_io_enable),
    .io_value(SaturatingCounter_271_io_value)
  );
  SaturatingCounter SaturatingCounter_272 (
    .clock(SaturatingCounter_272_clock),
    .reset(SaturatingCounter_272_reset),
    .io_enable(SaturatingCounter_272_io_enable),
    .io_value(SaturatingCounter_272_io_value)
  );
  SaturatingCounter SaturatingCounter_273 (
    .clock(SaturatingCounter_273_clock),
    .reset(SaturatingCounter_273_reset),
    .io_enable(SaturatingCounter_273_io_enable),
    .io_value(SaturatingCounter_273_io_value)
  );
  SaturatingCounter SaturatingCounter_274 (
    .clock(SaturatingCounter_274_clock),
    .reset(SaturatingCounter_274_reset),
    .io_enable(SaturatingCounter_274_io_enable),
    .io_value(SaturatingCounter_274_io_value)
  );
  SaturatingCounter SaturatingCounter_275 (
    .clock(SaturatingCounter_275_clock),
    .reset(SaturatingCounter_275_reset),
    .io_enable(SaturatingCounter_275_io_enable),
    .io_value(SaturatingCounter_275_io_value)
  );
  SaturatingCounter SaturatingCounter_276 (
    .clock(SaturatingCounter_276_clock),
    .reset(SaturatingCounter_276_reset),
    .io_enable(SaturatingCounter_276_io_enable),
    .io_value(SaturatingCounter_276_io_value)
  );
  SaturatingCounter SaturatingCounter_277 (
    .clock(SaturatingCounter_277_clock),
    .reset(SaturatingCounter_277_reset),
    .io_enable(SaturatingCounter_277_io_enable),
    .io_value(SaturatingCounter_277_io_value)
  );
  SaturatingCounter SaturatingCounter_278 (
    .clock(SaturatingCounter_278_clock),
    .reset(SaturatingCounter_278_reset),
    .io_enable(SaturatingCounter_278_io_enable),
    .io_value(SaturatingCounter_278_io_value)
  );
  SaturatingCounter SaturatingCounter_279 (
    .clock(SaturatingCounter_279_clock),
    .reset(SaturatingCounter_279_reset),
    .io_enable(SaturatingCounter_279_io_enable),
    .io_value(SaturatingCounter_279_io_value)
  );
  SaturatingCounter SaturatingCounter_280 (
    .clock(SaturatingCounter_280_clock),
    .reset(SaturatingCounter_280_reset),
    .io_enable(SaturatingCounter_280_io_enable),
    .io_value(SaturatingCounter_280_io_value)
  );
  SaturatingCounter SaturatingCounter_281 (
    .clock(SaturatingCounter_281_clock),
    .reset(SaturatingCounter_281_reset),
    .io_enable(SaturatingCounter_281_io_enable),
    .io_value(SaturatingCounter_281_io_value)
  );
  SaturatingCounter SaturatingCounter_282 (
    .clock(SaturatingCounter_282_clock),
    .reset(SaturatingCounter_282_reset),
    .io_enable(SaturatingCounter_282_io_enable),
    .io_value(SaturatingCounter_282_io_value)
  );
  SaturatingCounter SaturatingCounter_283 (
    .clock(SaturatingCounter_283_clock),
    .reset(SaturatingCounter_283_reset),
    .io_enable(SaturatingCounter_283_io_enable),
    .io_value(SaturatingCounter_283_io_value)
  );
  SaturatingCounter SaturatingCounter_284 (
    .clock(SaturatingCounter_284_clock),
    .reset(SaturatingCounter_284_reset),
    .io_enable(SaturatingCounter_284_io_enable),
    .io_value(SaturatingCounter_284_io_value)
  );
  SaturatingCounter SaturatingCounter_285 (
    .clock(SaturatingCounter_285_clock),
    .reset(SaturatingCounter_285_reset),
    .io_enable(SaturatingCounter_285_io_enable),
    .io_value(SaturatingCounter_285_io_value)
  );
  SaturatingCounter SaturatingCounter_286 (
    .clock(SaturatingCounter_286_clock),
    .reset(SaturatingCounter_286_reset),
    .io_enable(SaturatingCounter_286_io_enable),
    .io_value(SaturatingCounter_286_io_value)
  );
  SaturatingCounter SaturatingCounter_287 (
    .clock(SaturatingCounter_287_clock),
    .reset(SaturatingCounter_287_reset),
    .io_enable(SaturatingCounter_287_io_enable),
    .io_value(SaturatingCounter_287_io_value)
  );
  SaturatingCounter SaturatingCounter_288 (
    .clock(SaturatingCounter_288_clock),
    .reset(SaturatingCounter_288_reset),
    .io_enable(SaturatingCounter_288_io_enable),
    .io_value(SaturatingCounter_288_io_value)
  );
  SaturatingCounter SaturatingCounter_289 (
    .clock(SaturatingCounter_289_clock),
    .reset(SaturatingCounter_289_reset),
    .io_enable(SaturatingCounter_289_io_enable),
    .io_value(SaturatingCounter_289_io_value)
  );
  SaturatingCounter SaturatingCounter_290 (
    .clock(SaturatingCounter_290_clock),
    .reset(SaturatingCounter_290_reset),
    .io_enable(SaturatingCounter_290_io_enable),
    .io_value(SaturatingCounter_290_io_value)
  );
  SaturatingCounter SaturatingCounter_291 (
    .clock(SaturatingCounter_291_clock),
    .reset(SaturatingCounter_291_reset),
    .io_enable(SaturatingCounter_291_io_enable),
    .io_value(SaturatingCounter_291_io_value)
  );
  SaturatingCounter SaturatingCounter_292 (
    .clock(SaturatingCounter_292_clock),
    .reset(SaturatingCounter_292_reset),
    .io_enable(SaturatingCounter_292_io_enable),
    .io_value(SaturatingCounter_292_io_value)
  );
  SaturatingCounter SaturatingCounter_293 (
    .clock(SaturatingCounter_293_clock),
    .reset(SaturatingCounter_293_reset),
    .io_enable(SaturatingCounter_293_io_enable),
    .io_value(SaturatingCounter_293_io_value)
  );
  SaturatingCounter SaturatingCounter_294 (
    .clock(SaturatingCounter_294_clock),
    .reset(SaturatingCounter_294_reset),
    .io_enable(SaturatingCounter_294_io_enable),
    .io_value(SaturatingCounter_294_io_value)
  );
  SaturatingCounter SaturatingCounter_295 (
    .clock(SaturatingCounter_295_clock),
    .reset(SaturatingCounter_295_reset),
    .io_enable(SaturatingCounter_295_io_enable),
    .io_value(SaturatingCounter_295_io_value)
  );
  SaturatingCounter SaturatingCounter_296 (
    .clock(SaturatingCounter_296_clock),
    .reset(SaturatingCounter_296_reset),
    .io_enable(SaturatingCounter_296_io_enable),
    .io_value(SaturatingCounter_296_io_value)
  );
  SaturatingCounter SaturatingCounter_297 (
    .clock(SaturatingCounter_297_clock),
    .reset(SaturatingCounter_297_reset),
    .io_enable(SaturatingCounter_297_io_enable),
    .io_value(SaturatingCounter_297_io_value)
  );
  SaturatingCounter SaturatingCounter_298 (
    .clock(SaturatingCounter_298_clock),
    .reset(SaturatingCounter_298_reset),
    .io_enable(SaturatingCounter_298_io_enable),
    .io_value(SaturatingCounter_298_io_value)
  );
  SaturatingCounter SaturatingCounter_299 (
    .clock(SaturatingCounter_299_clock),
    .reset(SaturatingCounter_299_reset),
    .io_enable(SaturatingCounter_299_io_enable),
    .io_value(SaturatingCounter_299_io_value)
  );
  SaturatingCounter SaturatingCounter_300 (
    .clock(SaturatingCounter_300_clock),
    .reset(SaturatingCounter_300_reset),
    .io_enable(SaturatingCounter_300_io_enable),
    .io_value(SaturatingCounter_300_io_value)
  );
  SaturatingCounter SaturatingCounter_301 (
    .clock(SaturatingCounter_301_clock),
    .reset(SaturatingCounter_301_reset),
    .io_enable(SaturatingCounter_301_io_enable),
    .io_value(SaturatingCounter_301_io_value)
  );
  SaturatingCounter SaturatingCounter_302 (
    .clock(SaturatingCounter_302_clock),
    .reset(SaturatingCounter_302_reset),
    .io_enable(SaturatingCounter_302_io_enable),
    .io_value(SaturatingCounter_302_io_value)
  );
  SaturatingCounter SaturatingCounter_303 (
    .clock(SaturatingCounter_303_clock),
    .reset(SaturatingCounter_303_reset),
    .io_enable(SaturatingCounter_303_io_enable),
    .io_value(SaturatingCounter_303_io_value)
  );
  SaturatingCounter SaturatingCounter_304 (
    .clock(SaturatingCounter_304_clock),
    .reset(SaturatingCounter_304_reset),
    .io_enable(SaturatingCounter_304_io_enable),
    .io_value(SaturatingCounter_304_io_value)
  );
  SaturatingCounter SaturatingCounter_305 (
    .clock(SaturatingCounter_305_clock),
    .reset(SaturatingCounter_305_reset),
    .io_enable(SaturatingCounter_305_io_enable),
    .io_value(SaturatingCounter_305_io_value)
  );
  SaturatingCounter SaturatingCounter_306 (
    .clock(SaturatingCounter_306_clock),
    .reset(SaturatingCounter_306_reset),
    .io_enable(SaturatingCounter_306_io_enable),
    .io_value(SaturatingCounter_306_io_value)
  );
  SaturatingCounter SaturatingCounter_307 (
    .clock(SaturatingCounter_307_clock),
    .reset(SaturatingCounter_307_reset),
    .io_enable(SaturatingCounter_307_io_enable),
    .io_value(SaturatingCounter_307_io_value)
  );
  SaturatingCounter SaturatingCounter_308 (
    .clock(SaturatingCounter_308_clock),
    .reset(SaturatingCounter_308_reset),
    .io_enable(SaturatingCounter_308_io_enable),
    .io_value(SaturatingCounter_308_io_value)
  );
  SaturatingCounter SaturatingCounter_309 (
    .clock(SaturatingCounter_309_clock),
    .reset(SaturatingCounter_309_reset),
    .io_enable(SaturatingCounter_309_io_enable),
    .io_value(SaturatingCounter_309_io_value)
  );
  SaturatingCounter SaturatingCounter_310 (
    .clock(SaturatingCounter_310_clock),
    .reset(SaturatingCounter_310_reset),
    .io_enable(SaturatingCounter_310_io_enable),
    .io_value(SaturatingCounter_310_io_value)
  );
  SaturatingCounter SaturatingCounter_311 (
    .clock(SaturatingCounter_311_clock),
    .reset(SaturatingCounter_311_reset),
    .io_enable(SaturatingCounter_311_io_enable),
    .io_value(SaturatingCounter_311_io_value)
  );
  SaturatingCounter SaturatingCounter_312 (
    .clock(SaturatingCounter_312_clock),
    .reset(SaturatingCounter_312_reset),
    .io_enable(SaturatingCounter_312_io_enable),
    .io_value(SaturatingCounter_312_io_value)
  );
  SaturatingCounter SaturatingCounter_313 (
    .clock(SaturatingCounter_313_clock),
    .reset(SaturatingCounter_313_reset),
    .io_enable(SaturatingCounter_313_io_enable),
    .io_value(SaturatingCounter_313_io_value)
  );
  SaturatingCounter SaturatingCounter_314 (
    .clock(SaturatingCounter_314_clock),
    .reset(SaturatingCounter_314_reset),
    .io_enable(SaturatingCounter_314_io_enable),
    .io_value(SaturatingCounter_314_io_value)
  );
  SaturatingCounter SaturatingCounter_315 (
    .clock(SaturatingCounter_315_clock),
    .reset(SaturatingCounter_315_reset),
    .io_enable(SaturatingCounter_315_io_enable),
    .io_value(SaturatingCounter_315_io_value)
  );
  SaturatingCounter SaturatingCounter_316 (
    .clock(SaturatingCounter_316_clock),
    .reset(SaturatingCounter_316_reset),
    .io_enable(SaturatingCounter_316_io_enable),
    .io_value(SaturatingCounter_316_io_value)
  );
  SaturatingCounter SaturatingCounter_317 (
    .clock(SaturatingCounter_317_clock),
    .reset(SaturatingCounter_317_reset),
    .io_enable(SaturatingCounter_317_io_enable),
    .io_value(SaturatingCounter_317_io_value)
  );
  SaturatingCounter SaturatingCounter_318 (
    .clock(SaturatingCounter_318_clock),
    .reset(SaturatingCounter_318_reset),
    .io_enable(SaturatingCounter_318_io_enable),
    .io_value(SaturatingCounter_318_io_value)
  );
  SaturatingCounter SaturatingCounter_319 (
    .clock(SaturatingCounter_319_clock),
    .reset(SaturatingCounter_319_reset),
    .io_enable(SaturatingCounter_319_io_enable),
    .io_value(SaturatingCounter_319_io_value)
  );
  SaturatingCounter SaturatingCounter_320 (
    .clock(SaturatingCounter_320_clock),
    .reset(SaturatingCounter_320_reset),
    .io_enable(SaturatingCounter_320_io_enable),
    .io_value(SaturatingCounter_320_io_value)
  );
  SaturatingCounter SaturatingCounter_321 (
    .clock(SaturatingCounter_321_clock),
    .reset(SaturatingCounter_321_reset),
    .io_enable(SaturatingCounter_321_io_enable),
    .io_value(SaturatingCounter_321_io_value)
  );
  SaturatingCounter SaturatingCounter_322 (
    .clock(SaturatingCounter_322_clock),
    .reset(SaturatingCounter_322_reset),
    .io_enable(SaturatingCounter_322_io_enable),
    .io_value(SaturatingCounter_322_io_value)
  );
  SaturatingCounter SaturatingCounter_323 (
    .clock(SaturatingCounter_323_clock),
    .reset(SaturatingCounter_323_reset),
    .io_enable(SaturatingCounter_323_io_enable),
    .io_value(SaturatingCounter_323_io_value)
  );
  SaturatingCounter SaturatingCounter_324 (
    .clock(SaturatingCounter_324_clock),
    .reset(SaturatingCounter_324_reset),
    .io_enable(SaturatingCounter_324_io_enable),
    .io_value(SaturatingCounter_324_io_value)
  );
  SaturatingCounter SaturatingCounter_325 (
    .clock(SaturatingCounter_325_clock),
    .reset(SaturatingCounter_325_reset),
    .io_enable(SaturatingCounter_325_io_enable),
    .io_value(SaturatingCounter_325_io_value)
  );
  SaturatingCounter SaturatingCounter_326 (
    .clock(SaturatingCounter_326_clock),
    .reset(SaturatingCounter_326_reset),
    .io_enable(SaturatingCounter_326_io_enable),
    .io_value(SaturatingCounter_326_io_value)
  );
  SaturatingCounter SaturatingCounter_327 (
    .clock(SaturatingCounter_327_clock),
    .reset(SaturatingCounter_327_reset),
    .io_enable(SaturatingCounter_327_io_enable),
    .io_value(SaturatingCounter_327_io_value)
  );
  SaturatingCounter SaturatingCounter_328 (
    .clock(SaturatingCounter_328_clock),
    .reset(SaturatingCounter_328_reset),
    .io_enable(SaturatingCounter_328_io_enable),
    .io_value(SaturatingCounter_328_io_value)
  );
  SaturatingCounter SaturatingCounter_329 (
    .clock(SaturatingCounter_329_clock),
    .reset(SaturatingCounter_329_reset),
    .io_enable(SaturatingCounter_329_io_enable),
    .io_value(SaturatingCounter_329_io_value)
  );
  SaturatingCounter SaturatingCounter_330 (
    .clock(SaturatingCounter_330_clock),
    .reset(SaturatingCounter_330_reset),
    .io_enable(SaturatingCounter_330_io_enable),
    .io_value(SaturatingCounter_330_io_value)
  );
  SaturatingCounter SaturatingCounter_331 (
    .clock(SaturatingCounter_331_clock),
    .reset(SaturatingCounter_331_reset),
    .io_enable(SaturatingCounter_331_io_enable),
    .io_value(SaturatingCounter_331_io_value)
  );
  SaturatingCounter SaturatingCounter_332 (
    .clock(SaturatingCounter_332_clock),
    .reset(SaturatingCounter_332_reset),
    .io_enable(SaturatingCounter_332_io_enable),
    .io_value(SaturatingCounter_332_io_value)
  );
  SaturatingCounter SaturatingCounter_333 (
    .clock(SaturatingCounter_333_clock),
    .reset(SaturatingCounter_333_reset),
    .io_enable(SaturatingCounter_333_io_enable),
    .io_value(SaturatingCounter_333_io_value)
  );
  SaturatingCounter SaturatingCounter_334 (
    .clock(SaturatingCounter_334_clock),
    .reset(SaturatingCounter_334_reset),
    .io_enable(SaturatingCounter_334_io_enable),
    .io_value(SaturatingCounter_334_io_value)
  );
  SaturatingCounter SaturatingCounter_335 (
    .clock(SaturatingCounter_335_clock),
    .reset(SaturatingCounter_335_reset),
    .io_enable(SaturatingCounter_335_io_enable),
    .io_value(SaturatingCounter_335_io_value)
  );
  SaturatingCounter SaturatingCounter_336 (
    .clock(SaturatingCounter_336_clock),
    .reset(SaturatingCounter_336_reset),
    .io_enable(SaturatingCounter_336_io_enable),
    .io_value(SaturatingCounter_336_io_value)
  );
  SaturatingCounter SaturatingCounter_337 (
    .clock(SaturatingCounter_337_clock),
    .reset(SaturatingCounter_337_reset),
    .io_enable(SaturatingCounter_337_io_enable),
    .io_value(SaturatingCounter_337_io_value)
  );
  SaturatingCounter SaturatingCounter_338 (
    .clock(SaturatingCounter_338_clock),
    .reset(SaturatingCounter_338_reset),
    .io_enable(SaturatingCounter_338_io_enable),
    .io_value(SaturatingCounter_338_io_value)
  );
  SaturatingCounter SaturatingCounter_339 (
    .clock(SaturatingCounter_339_clock),
    .reset(SaturatingCounter_339_reset),
    .io_enable(SaturatingCounter_339_io_enable),
    .io_value(SaturatingCounter_339_io_value)
  );
  SaturatingCounter SaturatingCounter_340 (
    .clock(SaturatingCounter_340_clock),
    .reset(SaturatingCounter_340_reset),
    .io_enable(SaturatingCounter_340_io_enable),
    .io_value(SaturatingCounter_340_io_value)
  );
  SaturatingCounter SaturatingCounter_341 (
    .clock(SaturatingCounter_341_clock),
    .reset(SaturatingCounter_341_reset),
    .io_enable(SaturatingCounter_341_io_enable),
    .io_value(SaturatingCounter_341_io_value)
  );
  SaturatingCounter SaturatingCounter_342 (
    .clock(SaturatingCounter_342_clock),
    .reset(SaturatingCounter_342_reset),
    .io_enable(SaturatingCounter_342_io_enable),
    .io_value(SaturatingCounter_342_io_value)
  );
  SaturatingCounter SaturatingCounter_343 (
    .clock(SaturatingCounter_343_clock),
    .reset(SaturatingCounter_343_reset),
    .io_enable(SaturatingCounter_343_io_enable),
    .io_value(SaturatingCounter_343_io_value)
  );
  SaturatingCounter SaturatingCounter_344 (
    .clock(SaturatingCounter_344_clock),
    .reset(SaturatingCounter_344_reset),
    .io_enable(SaturatingCounter_344_io_enable),
    .io_value(SaturatingCounter_344_io_value)
  );
  SaturatingCounter SaturatingCounter_345 (
    .clock(SaturatingCounter_345_clock),
    .reset(SaturatingCounter_345_reset),
    .io_enable(SaturatingCounter_345_io_enable),
    .io_value(SaturatingCounter_345_io_value)
  );
  SaturatingCounter SaturatingCounter_346 (
    .clock(SaturatingCounter_346_clock),
    .reset(SaturatingCounter_346_reset),
    .io_enable(SaturatingCounter_346_io_enable),
    .io_value(SaturatingCounter_346_io_value)
  );
  SaturatingCounter SaturatingCounter_347 (
    .clock(SaturatingCounter_347_clock),
    .reset(SaturatingCounter_347_reset),
    .io_enable(SaturatingCounter_347_io_enable),
    .io_value(SaturatingCounter_347_io_value)
  );
  SaturatingCounter SaturatingCounter_348 (
    .clock(SaturatingCounter_348_clock),
    .reset(SaturatingCounter_348_reset),
    .io_enable(SaturatingCounter_348_io_enable),
    .io_value(SaturatingCounter_348_io_value)
  );
  SaturatingCounter SaturatingCounter_349 (
    .clock(SaturatingCounter_349_clock),
    .reset(SaturatingCounter_349_reset),
    .io_enable(SaturatingCounter_349_io_enable),
    .io_value(SaturatingCounter_349_io_value)
  );
  SaturatingCounter SaturatingCounter_350 (
    .clock(SaturatingCounter_350_clock),
    .reset(SaturatingCounter_350_reset),
    .io_enable(SaturatingCounter_350_io_enable),
    .io_value(SaturatingCounter_350_io_value)
  );
  SaturatingCounter SaturatingCounter_351 (
    .clock(SaturatingCounter_351_clock),
    .reset(SaturatingCounter_351_reset),
    .io_enable(SaturatingCounter_351_io_enable),
    .io_value(SaturatingCounter_351_io_value)
  );
  SaturatingCounter SaturatingCounter_352 (
    .clock(SaturatingCounter_352_clock),
    .reset(SaturatingCounter_352_reset),
    .io_enable(SaturatingCounter_352_io_enable),
    .io_value(SaturatingCounter_352_io_value)
  );
  SaturatingCounter SaturatingCounter_353 (
    .clock(SaturatingCounter_353_clock),
    .reset(SaturatingCounter_353_reset),
    .io_enable(SaturatingCounter_353_io_enable),
    .io_value(SaturatingCounter_353_io_value)
  );
  SaturatingCounter SaturatingCounter_354 (
    .clock(SaturatingCounter_354_clock),
    .reset(SaturatingCounter_354_reset),
    .io_enable(SaturatingCounter_354_io_enable),
    .io_value(SaturatingCounter_354_io_value)
  );
  SaturatingCounter SaturatingCounter_355 (
    .clock(SaturatingCounter_355_clock),
    .reset(SaturatingCounter_355_reset),
    .io_enable(SaturatingCounter_355_io_enable),
    .io_value(SaturatingCounter_355_io_value)
  );
  SaturatingCounter SaturatingCounter_356 (
    .clock(SaturatingCounter_356_clock),
    .reset(SaturatingCounter_356_reset),
    .io_enable(SaturatingCounter_356_io_enable),
    .io_value(SaturatingCounter_356_io_value)
  );
  SaturatingCounter SaturatingCounter_357 (
    .clock(SaturatingCounter_357_clock),
    .reset(SaturatingCounter_357_reset),
    .io_enable(SaturatingCounter_357_io_enable),
    .io_value(SaturatingCounter_357_io_value)
  );
  SaturatingCounter SaturatingCounter_358 (
    .clock(SaturatingCounter_358_clock),
    .reset(SaturatingCounter_358_reset),
    .io_enable(SaturatingCounter_358_io_enable),
    .io_value(SaturatingCounter_358_io_value)
  );
  SaturatingCounter SaturatingCounter_359 (
    .clock(SaturatingCounter_359_clock),
    .reset(SaturatingCounter_359_reset),
    .io_enable(SaturatingCounter_359_io_enable),
    .io_value(SaturatingCounter_359_io_value)
  );
  SaturatingCounter SaturatingCounter_360 (
    .clock(SaturatingCounter_360_clock),
    .reset(SaturatingCounter_360_reset),
    .io_enable(SaturatingCounter_360_io_enable),
    .io_value(SaturatingCounter_360_io_value)
  );
  SaturatingCounter SaturatingCounter_361 (
    .clock(SaturatingCounter_361_clock),
    .reset(SaturatingCounter_361_reset),
    .io_enable(SaturatingCounter_361_io_enable),
    .io_value(SaturatingCounter_361_io_value)
  );
  SaturatingCounter SaturatingCounter_362 (
    .clock(SaturatingCounter_362_clock),
    .reset(SaturatingCounter_362_reset),
    .io_enable(SaturatingCounter_362_io_enable),
    .io_value(SaturatingCounter_362_io_value)
  );
  SaturatingCounter SaturatingCounter_363 (
    .clock(SaturatingCounter_363_clock),
    .reset(SaturatingCounter_363_reset),
    .io_enable(SaturatingCounter_363_io_enable),
    .io_value(SaturatingCounter_363_io_value)
  );
  SaturatingCounter SaturatingCounter_364 (
    .clock(SaturatingCounter_364_clock),
    .reset(SaturatingCounter_364_reset),
    .io_enable(SaturatingCounter_364_io_enable),
    .io_value(SaturatingCounter_364_io_value)
  );
  SaturatingCounter SaturatingCounter_365 (
    .clock(SaturatingCounter_365_clock),
    .reset(SaturatingCounter_365_reset),
    .io_enable(SaturatingCounter_365_io_enable),
    .io_value(SaturatingCounter_365_io_value)
  );
  SaturatingCounter SaturatingCounter_366 (
    .clock(SaturatingCounter_366_clock),
    .reset(SaturatingCounter_366_reset),
    .io_enable(SaturatingCounter_366_io_enable),
    .io_value(SaturatingCounter_366_io_value)
  );
  SaturatingCounter SaturatingCounter_367 (
    .clock(SaturatingCounter_367_clock),
    .reset(SaturatingCounter_367_reset),
    .io_enable(SaturatingCounter_367_io_enable),
    .io_value(SaturatingCounter_367_io_value)
  );
  SaturatingCounter SaturatingCounter_368 (
    .clock(SaturatingCounter_368_clock),
    .reset(SaturatingCounter_368_reset),
    .io_enable(SaturatingCounter_368_io_enable),
    .io_value(SaturatingCounter_368_io_value)
  );
  SaturatingCounter SaturatingCounter_369 (
    .clock(SaturatingCounter_369_clock),
    .reset(SaturatingCounter_369_reset),
    .io_enable(SaturatingCounter_369_io_enable),
    .io_value(SaturatingCounter_369_io_value)
  );
  SaturatingCounter SaturatingCounter_370 (
    .clock(SaturatingCounter_370_clock),
    .reset(SaturatingCounter_370_reset),
    .io_enable(SaturatingCounter_370_io_enable),
    .io_value(SaturatingCounter_370_io_value)
  );
  SaturatingCounter SaturatingCounter_371 (
    .clock(SaturatingCounter_371_clock),
    .reset(SaturatingCounter_371_reset),
    .io_enable(SaturatingCounter_371_io_enable),
    .io_value(SaturatingCounter_371_io_value)
  );
  SaturatingCounter SaturatingCounter_372 (
    .clock(SaturatingCounter_372_clock),
    .reset(SaturatingCounter_372_reset),
    .io_enable(SaturatingCounter_372_io_enable),
    .io_value(SaturatingCounter_372_io_value)
  );
  SaturatingCounter SaturatingCounter_373 (
    .clock(SaturatingCounter_373_clock),
    .reset(SaturatingCounter_373_reset),
    .io_enable(SaturatingCounter_373_io_enable),
    .io_value(SaturatingCounter_373_io_value)
  );
  SaturatingCounter SaturatingCounter_374 (
    .clock(SaturatingCounter_374_clock),
    .reset(SaturatingCounter_374_reset),
    .io_enable(SaturatingCounter_374_io_enable),
    .io_value(SaturatingCounter_374_io_value)
  );
  SaturatingCounter SaturatingCounter_375 (
    .clock(SaturatingCounter_375_clock),
    .reset(SaturatingCounter_375_reset),
    .io_enable(SaturatingCounter_375_io_enable),
    .io_value(SaturatingCounter_375_io_value)
  );
  SaturatingCounter SaturatingCounter_376 (
    .clock(SaturatingCounter_376_clock),
    .reset(SaturatingCounter_376_reset),
    .io_enable(SaturatingCounter_376_io_enable),
    .io_value(SaturatingCounter_376_io_value)
  );
  SaturatingCounter SaturatingCounter_377 (
    .clock(SaturatingCounter_377_clock),
    .reset(SaturatingCounter_377_reset),
    .io_enable(SaturatingCounter_377_io_enable),
    .io_value(SaturatingCounter_377_io_value)
  );
  SaturatingCounter SaturatingCounter_378 (
    .clock(SaturatingCounter_378_clock),
    .reset(SaturatingCounter_378_reset),
    .io_enable(SaturatingCounter_378_io_enable),
    .io_value(SaturatingCounter_378_io_value)
  );
  SaturatingCounter SaturatingCounter_379 (
    .clock(SaturatingCounter_379_clock),
    .reset(SaturatingCounter_379_reset),
    .io_enable(SaturatingCounter_379_io_enable),
    .io_value(SaturatingCounter_379_io_value)
  );
  SaturatingCounter SaturatingCounter_380 (
    .clock(SaturatingCounter_380_clock),
    .reset(SaturatingCounter_380_reset),
    .io_enable(SaturatingCounter_380_io_enable),
    .io_value(SaturatingCounter_380_io_value)
  );
  SaturatingCounter SaturatingCounter_381 (
    .clock(SaturatingCounter_381_clock),
    .reset(SaturatingCounter_381_reset),
    .io_enable(SaturatingCounter_381_io_enable),
    .io_value(SaturatingCounter_381_io_value)
  );
  SaturatingCounter SaturatingCounter_382 (
    .clock(SaturatingCounter_382_clock),
    .reset(SaturatingCounter_382_reset),
    .io_enable(SaturatingCounter_382_io_enable),
    .io_value(SaturatingCounter_382_io_value)
  );
  assign _T_219 = {io_input_bytes_6,io_input_bytes_7};
  assign _T_220 = {io_input_bytes_4,io_input_bytes_5};
  assign _T_221 = {_T_220,_T_219};
  assign _T_222 = {io_input_bytes_2,io_input_bytes_3};
  assign _T_223 = {io_input_bytes_0,io_input_bytes_1};
  assign _T_224 = {_T_223,_T_222};
  assign input_bytes = {_T_224,_T_221};
  assign _T_225 = input_bytes[63:29];
  assign _T_227 = dut_io_coverage_0;
  assign coverage_0 = {7'h0,SaturatingCounter_io_value};
  assign _T_232 = dut_io_coverage_1;
  assign _T_233 = ~ dut_io_coverage_1;
  assign _T_237 = {6'h0,SaturatingCounter_1_io_value};
  assign coverage_1 = {_T_237,SaturatingCounter_2_io_value};
  assign _T_239 = dut_io_coverage_2;
  assign _T_240 = ~ dut_io_coverage_2;
  assign _T_244 = {6'h0,SaturatingCounter_3_io_value};
  assign coverage_2 = {_T_244,SaturatingCounter_4_io_value};
  assign _T_246 = dut_io_coverage_3;
  assign _T_247 = ~ dut_io_coverage_3;
  assign _T_251 = {6'h0,SaturatingCounter_5_io_value};
  assign coverage_3 = {_T_251,SaturatingCounter_6_io_value};
  assign _T_253 = dut_io_coverage_4;
  assign _T_254 = ~ dut_io_coverage_4;
  assign _T_258 = {6'h0,SaturatingCounter_7_io_value};
  assign coverage_4 = {_T_258,SaturatingCounter_8_io_value};
  assign _T_260 = dut_io_coverage_5;
  assign _T_261 = ~ dut_io_coverage_5;
  assign _T_265 = {6'h0,SaturatingCounter_9_io_value};
  assign coverage_5 = {_T_265,SaturatingCounter_10_io_value};
  assign _T_267 = dut_io_coverage_6;
  assign _T_268 = ~ dut_io_coverage_6;
  assign _T_272 = {6'h0,SaturatingCounter_11_io_value};
  assign coverage_6 = {_T_272,SaturatingCounter_12_io_value};
  assign _T_274 = dut_io_coverage_7;
  assign _T_275 = ~ dut_io_coverage_7;
  assign _T_279 = {6'h0,SaturatingCounter_13_io_value};
  assign coverage_7 = {_T_279,SaturatingCounter_14_io_value};
  assign _T_281 = dut_io_coverage_8;
  assign _T_282 = ~ dut_io_coverage_8;
  assign _T_286 = {6'h0,SaturatingCounter_15_io_value};
  assign coverage_8 = {_T_286,SaturatingCounter_16_io_value};
  assign _T_288 = dut_io_coverage_9;
  assign _T_289 = ~ dut_io_coverage_9;
  assign _T_293 = {6'h0,SaturatingCounter_17_io_value};
  assign coverage_9 = {_T_293,SaturatingCounter_18_io_value};
  assign _T_295 = dut_io_coverage_10;
  assign _T_296 = ~ dut_io_coverage_10;
  assign _T_300 = {6'h0,SaturatingCounter_19_io_value};
  assign coverage_10 = {_T_300,SaturatingCounter_20_io_value};
  assign _T_302 = dut_io_coverage_11;
  assign _T_303 = ~ dut_io_coverage_11;
  assign _T_307 = {6'h0,SaturatingCounter_21_io_value};
  assign coverage_11 = {_T_307,SaturatingCounter_22_io_value};
  assign _T_309 = dut_io_coverage_12;
  assign _T_310 = ~ dut_io_coverage_12;
  assign _T_314 = {6'h0,SaturatingCounter_23_io_value};
  assign coverage_12 = {_T_314,SaturatingCounter_24_io_value};
  assign _T_316 = dut_io_coverage_13;
  assign _T_317 = ~ dut_io_coverage_13;
  assign _T_321 = {6'h0,SaturatingCounter_25_io_value};
  assign coverage_13 = {_T_321,SaturatingCounter_26_io_value};
  assign _T_323 = dut_io_coverage_14;
  assign _T_324 = ~ dut_io_coverage_14;
  assign _T_328 = {6'h0,SaturatingCounter_27_io_value};
  assign coverage_14 = {_T_328,SaturatingCounter_28_io_value};
  assign _T_330 = dut_io_coverage_15;
  assign _T_331 = ~ dut_io_coverage_15;
  assign _T_335 = {6'h0,SaturatingCounter_29_io_value};
  assign coverage_15 = {_T_335,SaturatingCounter_30_io_value};
  assign _T_337 = dut_io_coverage_16;
  assign _T_338 = ~ dut_io_coverage_16;
  assign _T_342 = {6'h0,SaturatingCounter_31_io_value};
  assign coverage_16 = {_T_342,SaturatingCounter_32_io_value};
  assign _T_344 = dut_io_coverage_17;
  assign _T_345 = ~ dut_io_coverage_17;
  assign _T_349 = {6'h0,SaturatingCounter_33_io_value};
  assign coverage_17 = {_T_349,SaturatingCounter_34_io_value};
  assign _T_351 = dut_io_coverage_18;
  assign _T_352 = ~ dut_io_coverage_18;
  assign _T_356 = {6'h0,SaturatingCounter_35_io_value};
  assign coverage_18 = {_T_356,SaturatingCounter_36_io_value};
  assign _T_358 = dut_io_coverage_19;
  assign _T_359 = ~ dut_io_coverage_19;
  assign _T_363 = {6'h0,SaturatingCounter_37_io_value};
  assign coverage_19 = {_T_363,SaturatingCounter_38_io_value};
  assign _T_365 = dut_io_coverage_20;
  assign _T_366 = ~ dut_io_coverage_20;
  assign _T_370 = {6'h0,SaturatingCounter_39_io_value};
  assign coverage_20 = {_T_370,SaturatingCounter_40_io_value};
  assign _T_372 = dut_io_coverage_21;
  assign _T_373 = ~ dut_io_coverage_21;
  assign _T_377 = {6'h0,SaturatingCounter_41_io_value};
  assign coverage_21 = {_T_377,SaturatingCounter_42_io_value};
  assign _T_379 = dut_io_coverage_22;
  assign _T_380 = ~ dut_io_coverage_22;
  assign _T_384 = {6'h0,SaturatingCounter_43_io_value};
  assign coverage_22 = {_T_384,SaturatingCounter_44_io_value};
  assign _T_386 = dut_io_coverage_23;
  assign _T_387 = ~ dut_io_coverage_23;
  assign _T_391 = {6'h0,SaturatingCounter_45_io_value};
  assign coverage_23 = {_T_391,SaturatingCounter_46_io_value};
  assign _T_393 = dut_io_coverage_24;
  assign _T_394 = ~ dut_io_coverage_24;
  assign _T_398 = {6'h0,SaturatingCounter_47_io_value};
  assign coverage_24 = {_T_398,SaturatingCounter_48_io_value};
  assign _T_400 = dut_io_coverage_25;
  assign _T_401 = ~ dut_io_coverage_25;
  assign _T_405 = {6'h0,SaturatingCounter_49_io_value};
  assign coverage_25 = {_T_405,SaturatingCounter_50_io_value};
  assign _T_407 = dut_io_coverage_26;
  assign _T_408 = ~ dut_io_coverage_26;
  assign _T_412 = {6'h0,SaturatingCounter_51_io_value};
  assign coverage_26 = {_T_412,SaturatingCounter_52_io_value};
  assign _T_414 = dut_io_coverage_27;
  assign _T_415 = ~ dut_io_coverage_27;
  assign _T_419 = {6'h0,SaturatingCounter_53_io_value};
  assign coverage_27 = {_T_419,SaturatingCounter_54_io_value};
  assign _T_421 = dut_io_coverage_28;
  assign _T_422 = ~ dut_io_coverage_28;
  assign _T_426 = {6'h0,SaturatingCounter_55_io_value};
  assign coverage_28 = {_T_426,SaturatingCounter_56_io_value};
  assign _T_428 = dut_io_coverage_29;
  assign _T_429 = ~ dut_io_coverage_29;
  assign _T_433 = {6'h0,SaturatingCounter_57_io_value};
  assign coverage_29 = {_T_433,SaturatingCounter_58_io_value};
  assign _T_435 = dut_io_coverage_30;
  assign _T_436 = ~ dut_io_coverage_30;
  assign _T_440 = {6'h0,SaturatingCounter_59_io_value};
  assign coverage_30 = {_T_440,SaturatingCounter_60_io_value};
  assign _T_442 = dut_io_coverage_31;
  assign _T_443 = ~ dut_io_coverage_31;
  assign _T_447 = {6'h0,SaturatingCounter_61_io_value};
  assign coverage_31 = {_T_447,SaturatingCounter_62_io_value};
  assign _T_449 = dut_io_coverage_32;
  assign _T_450 = ~ dut_io_coverage_32;
  assign _T_454 = {6'h0,SaturatingCounter_63_io_value};
  assign coverage_32 = {_T_454,SaturatingCounter_64_io_value};
  assign _T_456 = dut_io_coverage_33;
  assign _T_457 = ~ dut_io_coverage_33;
  assign _T_461 = {6'h0,SaturatingCounter_65_io_value};
  assign coverage_33 = {_T_461,SaturatingCounter_66_io_value};
  assign _T_463 = dut_io_coverage_34;
  assign _T_464 = ~ dut_io_coverage_34;
  assign _T_468 = {6'h0,SaturatingCounter_67_io_value};
  assign coverage_34 = {_T_468,SaturatingCounter_68_io_value};
  assign _T_470 = dut_io_coverage_35;
  assign _T_471 = ~ dut_io_coverage_35;
  assign _T_475 = {6'h0,SaturatingCounter_69_io_value};
  assign coverage_35 = {_T_475,SaturatingCounter_70_io_value};
  assign _T_477 = dut_io_coverage_36;
  assign _T_478 = ~ dut_io_coverage_36;
  assign _T_482 = {6'h0,SaturatingCounter_71_io_value};
  assign coverage_36 = {_T_482,SaturatingCounter_72_io_value};
  assign _T_484 = dut_io_coverage_37;
  assign _T_485 = ~ dut_io_coverage_37;
  assign _T_489 = {6'h0,SaturatingCounter_73_io_value};
  assign coverage_37 = {_T_489,SaturatingCounter_74_io_value};
  assign _T_491 = dut_io_coverage_38;
  assign _T_492 = ~ dut_io_coverage_38;
  assign _T_496 = {6'h0,SaturatingCounter_75_io_value};
  assign coverage_38 = {_T_496,SaturatingCounter_76_io_value};
  assign _T_498 = dut_io_coverage_39;
  assign _T_499 = ~ dut_io_coverage_39;
  assign _T_503 = {6'h0,SaturatingCounter_77_io_value};
  assign coverage_39 = {_T_503,SaturatingCounter_78_io_value};
  assign _T_505 = dut_io_coverage_40;
  assign _T_506 = ~ dut_io_coverage_40;
  assign _T_510 = {6'h0,SaturatingCounter_79_io_value};
  assign coverage_40 = {_T_510,SaturatingCounter_80_io_value};
  assign _T_512 = dut_io_coverage_41;
  assign _T_513 = ~ dut_io_coverage_41;
  assign _T_517 = {6'h0,SaturatingCounter_81_io_value};
  assign coverage_41 = {_T_517,SaturatingCounter_82_io_value};
  assign _T_519 = dut_io_coverage_42;
  assign _T_520 = ~ dut_io_coverage_42;
  assign _T_524 = {6'h0,SaturatingCounter_83_io_value};
  assign coverage_42 = {_T_524,SaturatingCounter_84_io_value};
  assign _T_526 = dut_io_coverage_43;
  assign _T_527 = ~ dut_io_coverage_43;
  assign _T_531 = {6'h0,SaturatingCounter_85_io_value};
  assign coverage_43 = {_T_531,SaturatingCounter_86_io_value};
  assign _T_533 = dut_io_coverage_44;
  assign _T_534 = ~ dut_io_coverage_44;
  assign _T_538 = {6'h0,SaturatingCounter_87_io_value};
  assign coverage_44 = {_T_538,SaturatingCounter_88_io_value};
  assign _T_540 = dut_io_coverage_45;
  assign _T_541 = ~ dut_io_coverage_45;
  assign _T_545 = {6'h0,SaturatingCounter_89_io_value};
  assign coverage_45 = {_T_545,SaturatingCounter_90_io_value};
  assign _T_547 = dut_io_coverage_46;
  assign _T_548 = ~ dut_io_coverage_46;
  assign _T_552 = {6'h0,SaturatingCounter_91_io_value};
  assign coverage_46 = {_T_552,SaturatingCounter_92_io_value};
  assign _T_554 = dut_io_coverage_47;
  assign _T_555 = ~ dut_io_coverage_47;
  assign _T_559 = {6'h0,SaturatingCounter_93_io_value};
  assign coverage_47 = {_T_559,SaturatingCounter_94_io_value};
  assign _T_561 = dut_io_coverage_48;
  assign _T_562 = ~ dut_io_coverage_48;
  assign _T_566 = {6'h0,SaturatingCounter_95_io_value};
  assign coverage_48 = {_T_566,SaturatingCounter_96_io_value};
  assign _T_568 = dut_io_coverage_49;
  assign _T_569 = ~ dut_io_coverage_49;
  assign _T_573 = {6'h0,SaturatingCounter_97_io_value};
  assign coverage_49 = {_T_573,SaturatingCounter_98_io_value};
  assign _T_575 = dut_io_coverage_50;
  assign _T_576 = ~ dut_io_coverage_50;
  assign _T_580 = {6'h0,SaturatingCounter_99_io_value};
  assign coverage_50 = {_T_580,SaturatingCounter_100_io_value};
  assign _T_582 = dut_io_coverage_51;
  assign _T_583 = ~ dut_io_coverage_51;
  assign _T_587 = {6'h0,SaturatingCounter_101_io_value};
  assign coverage_51 = {_T_587,SaturatingCounter_102_io_value};
  assign _T_589 = dut_io_coverage_52;
  assign _T_590 = ~ dut_io_coverage_52;
  assign _T_594 = {6'h0,SaturatingCounter_103_io_value};
  assign coverage_52 = {_T_594,SaturatingCounter_104_io_value};
  assign _T_596 = dut_io_coverage_53;
  assign _T_597 = ~ dut_io_coverage_53;
  assign _T_601 = {6'h0,SaturatingCounter_105_io_value};
  assign coverage_53 = {_T_601,SaturatingCounter_106_io_value};
  assign _T_603 = dut_io_coverage_54;
  assign _T_604 = ~ dut_io_coverage_54;
  assign _T_608 = {6'h0,SaturatingCounter_107_io_value};
  assign coverage_54 = {_T_608,SaturatingCounter_108_io_value};
  assign _T_610 = dut_io_coverage_55;
  assign _T_611 = ~ dut_io_coverage_55;
  assign _T_615 = {6'h0,SaturatingCounter_109_io_value};
  assign coverage_55 = {_T_615,SaturatingCounter_110_io_value};
  assign _T_617 = dut_io_coverage_56;
  assign _T_618 = ~ dut_io_coverage_56;
  assign _T_622 = {6'h0,SaturatingCounter_111_io_value};
  assign coverage_56 = {_T_622,SaturatingCounter_112_io_value};
  assign _T_624 = dut_io_coverage_57;
  assign _T_625 = ~ dut_io_coverage_57;
  assign _T_629 = {6'h0,SaturatingCounter_113_io_value};
  assign coverage_57 = {_T_629,SaturatingCounter_114_io_value};
  assign _T_631 = dut_io_coverage_58;
  assign _T_632 = ~ dut_io_coverage_58;
  assign _T_636 = {6'h0,SaturatingCounter_115_io_value};
  assign coverage_58 = {_T_636,SaturatingCounter_116_io_value};
  assign _T_638 = dut_io_coverage_59;
  assign _T_639 = ~ dut_io_coverage_59;
  assign _T_643 = {6'h0,SaturatingCounter_117_io_value};
  assign coverage_59 = {_T_643,SaturatingCounter_118_io_value};
  assign _T_645 = dut_io_coverage_60;
  assign _T_646 = ~ dut_io_coverage_60;
  assign _T_650 = {6'h0,SaturatingCounter_119_io_value};
  assign coverage_60 = {_T_650,SaturatingCounter_120_io_value};
  assign _T_652 = dut_io_coverage_61;
  assign _T_653 = ~ dut_io_coverage_61;
  assign _T_657 = {6'h0,SaturatingCounter_121_io_value};
  assign coverage_61 = {_T_657,SaturatingCounter_122_io_value};
  assign _T_659 = dut_io_coverage_62;
  assign _T_660 = ~ dut_io_coverage_62;
  assign _T_664 = {6'h0,SaturatingCounter_123_io_value};
  assign coverage_62 = {_T_664,SaturatingCounter_124_io_value};
  assign _T_666 = dut_io_coverage_63;
  assign _T_667 = ~ dut_io_coverage_63;
  assign _T_671 = {6'h0,SaturatingCounter_125_io_value};
  assign coverage_63 = {_T_671,SaturatingCounter_126_io_value};
  assign _T_673 = dut_io_coverage_64;
  assign _T_674 = ~ dut_io_coverage_64;
  assign _T_678 = {6'h0,SaturatingCounter_127_io_value};
  assign coverage_64 = {_T_678,SaturatingCounter_128_io_value};
  assign _T_680 = dut_io_coverage_65;
  assign _T_681 = ~ dut_io_coverage_65;
  assign _T_685 = {6'h0,SaturatingCounter_129_io_value};
  assign coverage_65 = {_T_685,SaturatingCounter_130_io_value};
  assign _T_687 = dut_io_coverage_66;
  assign _T_688 = ~ dut_io_coverage_66;
  assign _T_692 = {6'h0,SaturatingCounter_131_io_value};
  assign coverage_66 = {_T_692,SaturatingCounter_132_io_value};
  assign _T_694 = dut_io_coverage_67;
  assign _T_695 = ~ dut_io_coverage_67;
  assign _T_699 = {6'h0,SaturatingCounter_133_io_value};
  assign coverage_67 = {_T_699,SaturatingCounter_134_io_value};
  assign _T_701 = dut_io_coverage_68;
  assign _T_702 = ~ dut_io_coverage_68;
  assign _T_706 = {6'h0,SaturatingCounter_135_io_value};
  assign coverage_68 = {_T_706,SaturatingCounter_136_io_value};
  assign _T_708 = dut_io_coverage_69;
  assign _T_709 = ~ dut_io_coverage_69;
  assign _T_713 = {6'h0,SaturatingCounter_137_io_value};
  assign coverage_69 = {_T_713,SaturatingCounter_138_io_value};
  assign _T_715 = dut_io_coverage_70;
  assign _T_716 = ~ dut_io_coverage_70;
  assign _T_720 = {6'h0,SaturatingCounter_139_io_value};
  assign coverage_70 = {_T_720,SaturatingCounter_140_io_value};
  assign _T_722 = dut_io_coverage_71;
  assign _T_723 = ~ dut_io_coverage_71;
  assign _T_727 = {6'h0,SaturatingCounter_141_io_value};
  assign coverage_71 = {_T_727,SaturatingCounter_142_io_value};
  assign _T_729 = dut_io_coverage_72;
  assign _T_730 = ~ dut_io_coverage_72;
  assign _T_734 = {6'h0,SaturatingCounter_143_io_value};
  assign coverage_72 = {_T_734,SaturatingCounter_144_io_value};
  assign _T_736 = dut_io_coverage_73;
  assign _T_737 = ~ dut_io_coverage_73;
  assign _T_741 = {6'h0,SaturatingCounter_145_io_value};
  assign coverage_73 = {_T_741,SaturatingCounter_146_io_value};
  assign _T_743 = dut_io_coverage_74;
  assign _T_744 = ~ dut_io_coverage_74;
  assign _T_748 = {6'h0,SaturatingCounter_147_io_value};
  assign coverage_74 = {_T_748,SaturatingCounter_148_io_value};
  assign _T_750 = dut_io_coverage_75;
  assign _T_751 = ~ dut_io_coverage_75;
  assign _T_755 = {6'h0,SaturatingCounter_149_io_value};
  assign coverage_75 = {_T_755,SaturatingCounter_150_io_value};
  assign _T_757 = dut_io_coverage_76;
  assign _T_758 = ~ dut_io_coverage_76;
  assign _T_762 = {6'h0,SaturatingCounter_151_io_value};
  assign coverage_76 = {_T_762,SaturatingCounter_152_io_value};
  assign _T_764 = dut_io_coverage_77;
  assign _T_765 = ~ dut_io_coverage_77;
  assign _T_769 = {6'h0,SaturatingCounter_153_io_value};
  assign coverage_77 = {_T_769,SaturatingCounter_154_io_value};
  assign _T_771 = dut_io_coverage_78;
  assign _T_772 = ~ dut_io_coverage_78;
  assign _T_776 = {6'h0,SaturatingCounter_155_io_value};
  assign coverage_78 = {_T_776,SaturatingCounter_156_io_value};
  assign _T_778 = dut_io_coverage_79;
  assign _T_779 = ~ dut_io_coverage_79;
  assign _T_783 = {6'h0,SaturatingCounter_157_io_value};
  assign coverage_79 = {_T_783,SaturatingCounter_158_io_value};
  assign _T_785 = dut_io_coverage_80;
  assign _T_786 = ~ dut_io_coverage_80;
  assign _T_790 = {6'h0,SaturatingCounter_159_io_value};
  assign coverage_80 = {_T_790,SaturatingCounter_160_io_value};
  assign _T_792 = dut_io_coverage_81;
  assign _T_793 = ~ dut_io_coverage_81;
  assign _T_797 = {6'h0,SaturatingCounter_161_io_value};
  assign coverage_81 = {_T_797,SaturatingCounter_162_io_value};
  assign _T_799 = dut_io_coverage_82;
  assign _T_800 = ~ dut_io_coverage_82;
  assign _T_804 = {6'h0,SaturatingCounter_163_io_value};
  assign coverage_82 = {_T_804,SaturatingCounter_164_io_value};
  assign _T_806 = dut_io_coverage_83;
  assign _T_807 = ~ dut_io_coverage_83;
  assign _T_811 = {6'h0,SaturatingCounter_165_io_value};
  assign coverage_83 = {_T_811,SaturatingCounter_166_io_value};
  assign _T_813 = dut_io_coverage_84;
  assign _T_814 = ~ dut_io_coverage_84;
  assign _T_818 = {6'h0,SaturatingCounter_167_io_value};
  assign coverage_84 = {_T_818,SaturatingCounter_168_io_value};
  assign _T_820 = dut_io_coverage_85;
  assign _T_821 = ~ dut_io_coverage_85;
  assign _T_825 = {6'h0,SaturatingCounter_169_io_value};
  assign coverage_85 = {_T_825,SaturatingCounter_170_io_value};
  assign _T_827 = dut_io_coverage_86;
  assign _T_828 = ~ dut_io_coverage_86;
  assign _T_832 = {6'h0,SaturatingCounter_171_io_value};
  assign coverage_86 = {_T_832,SaturatingCounter_172_io_value};
  assign _T_834 = dut_io_coverage_87;
  assign _T_835 = ~ dut_io_coverage_87;
  assign _T_839 = {6'h0,SaturatingCounter_173_io_value};
  assign coverage_87 = {_T_839,SaturatingCounter_174_io_value};
  assign _T_841 = dut_io_coverage_88;
  assign _T_842 = ~ dut_io_coverage_88;
  assign _T_846 = {6'h0,SaturatingCounter_175_io_value};
  assign coverage_88 = {_T_846,SaturatingCounter_176_io_value};
  assign _T_848 = dut_io_coverage_89;
  assign _T_849 = ~ dut_io_coverage_89;
  assign _T_853 = {6'h0,SaturatingCounter_177_io_value};
  assign coverage_89 = {_T_853,SaturatingCounter_178_io_value};
  assign _T_855 = dut_io_coverage_90;
  assign _T_856 = ~ dut_io_coverage_90;
  assign _T_860 = {6'h0,SaturatingCounter_179_io_value};
  assign coverage_90 = {_T_860,SaturatingCounter_180_io_value};
  assign _T_862 = dut_io_coverage_91;
  assign _T_863 = ~ dut_io_coverage_91;
  assign _T_867 = {6'h0,SaturatingCounter_181_io_value};
  assign coverage_91 = {_T_867,SaturatingCounter_182_io_value};
  assign _T_869 = dut_io_coverage_92;
  assign _T_870 = ~ dut_io_coverage_92;
  assign _T_874 = {6'h0,SaturatingCounter_183_io_value};
  assign coverage_92 = {_T_874,SaturatingCounter_184_io_value};
  assign _T_876 = dut_io_coverage_93;
  assign _T_877 = ~ dut_io_coverage_93;
  assign _T_881 = {6'h0,SaturatingCounter_185_io_value};
  assign coverage_93 = {_T_881,SaturatingCounter_186_io_value};
  assign _T_883 = dut_io_coverage_94;
  assign _T_884 = ~ dut_io_coverage_94;
  assign _T_888 = {6'h0,SaturatingCounter_187_io_value};
  assign coverage_94 = {_T_888,SaturatingCounter_188_io_value};
  assign _T_890 = dut_io_coverage_95;
  assign _T_891 = ~ dut_io_coverage_95;
  assign _T_895 = {6'h0,SaturatingCounter_189_io_value};
  assign coverage_95 = {_T_895,SaturatingCounter_190_io_value};
  assign _T_897 = dut_io_coverage_96;
  assign _T_898 = ~ dut_io_coverage_96;
  assign _T_902 = {6'h0,SaturatingCounter_191_io_value};
  assign coverage_96 = {_T_902,SaturatingCounter_192_io_value};
  assign _T_904 = dut_io_coverage_97;
  assign _T_905 = ~ dut_io_coverage_97;
  assign _T_909 = {6'h0,SaturatingCounter_193_io_value};
  assign coverage_97 = {_T_909,SaturatingCounter_194_io_value};
  assign _T_911 = dut_io_coverage_98;
  assign _T_912 = ~ dut_io_coverage_98;
  assign _T_916 = {6'h0,SaturatingCounter_195_io_value};
  assign coverage_98 = {_T_916,SaturatingCounter_196_io_value};
  assign _T_918 = dut_io_coverage_99;
  assign _T_919 = ~ dut_io_coverage_99;
  assign _T_923 = {6'h0,SaturatingCounter_197_io_value};
  assign coverage_99 = {_T_923,SaturatingCounter_198_io_value};
  assign _T_925 = dut_io_coverage_100;
  assign _T_926 = ~ dut_io_coverage_100;
  assign _T_930 = {6'h0,SaturatingCounter_199_io_value};
  assign coverage_100 = {_T_930,SaturatingCounter_200_io_value};
  assign _T_932 = dut_io_coverage_101;
  assign _T_933 = ~ dut_io_coverage_101;
  assign _T_937 = {6'h0,SaturatingCounter_201_io_value};
  assign coverage_101 = {_T_937,SaturatingCounter_202_io_value};
  assign _T_939 = dut_io_coverage_102;
  assign _T_940 = ~ dut_io_coverage_102;
  assign _T_944 = {6'h0,SaturatingCounter_203_io_value};
  assign coverage_102 = {_T_944,SaturatingCounter_204_io_value};
  assign _T_946 = dut_io_coverage_103;
  assign _T_947 = ~ dut_io_coverage_103;
  assign _T_951 = {6'h0,SaturatingCounter_205_io_value};
  assign coverage_103 = {_T_951,SaturatingCounter_206_io_value};
  assign _T_953 = dut_io_coverage_104;
  assign _T_954 = ~ dut_io_coverage_104;
  assign _T_958 = {6'h0,SaturatingCounter_207_io_value};
  assign coverage_104 = {_T_958,SaturatingCounter_208_io_value};
  assign _T_960 = dut_io_coverage_105;
  assign _T_961 = ~ dut_io_coverage_105;
  assign _T_965 = {6'h0,SaturatingCounter_209_io_value};
  assign coverage_105 = {_T_965,SaturatingCounter_210_io_value};
  assign _T_967 = dut_io_coverage_106;
  assign _T_968 = ~ dut_io_coverage_106;
  assign _T_972 = {6'h0,SaturatingCounter_211_io_value};
  assign coverage_106 = {_T_972,SaturatingCounter_212_io_value};
  assign _T_974 = dut_io_coverage_107;
  assign _T_975 = ~ dut_io_coverage_107;
  assign _T_979 = {6'h0,SaturatingCounter_213_io_value};
  assign coverage_107 = {_T_979,SaturatingCounter_214_io_value};
  assign _T_981 = dut_io_coverage_108;
  assign _T_982 = ~ dut_io_coverage_108;
  assign _T_986 = {6'h0,SaturatingCounter_215_io_value};
  assign coverage_108 = {_T_986,SaturatingCounter_216_io_value};
  assign _T_988 = dut_io_coverage_109;
  assign _T_989 = ~ dut_io_coverage_109;
  assign _T_993 = {6'h0,SaturatingCounter_217_io_value};
  assign coverage_109 = {_T_993,SaturatingCounter_218_io_value};
  assign _T_995 = dut_io_coverage_110;
  assign _T_996 = ~ dut_io_coverage_110;
  assign _T_1000 = {6'h0,SaturatingCounter_219_io_value};
  assign coverage_110 = {_T_1000,SaturatingCounter_220_io_value};
  assign _T_1002 = dut_io_coverage_111;
  assign _T_1003 = ~ dut_io_coverage_111;
  assign _T_1007 = {6'h0,SaturatingCounter_221_io_value};
  assign coverage_111 = {_T_1007,SaturatingCounter_222_io_value};
  assign _T_1009 = dut_io_coverage_112;
  assign _T_1010 = ~ dut_io_coverage_112;
  assign _T_1014 = {6'h0,SaturatingCounter_223_io_value};
  assign coverage_112 = {_T_1014,SaturatingCounter_224_io_value};
  assign _T_1016 = dut_io_coverage_113;
  assign _T_1017 = ~ dut_io_coverage_113;
  assign _T_1021 = {6'h0,SaturatingCounter_225_io_value};
  assign coverage_113 = {_T_1021,SaturatingCounter_226_io_value};
  assign _T_1023 = dut_io_coverage_114;
  assign _T_1024 = ~ dut_io_coverage_114;
  assign _T_1028 = {6'h0,SaturatingCounter_227_io_value};
  assign coverage_114 = {_T_1028,SaturatingCounter_228_io_value};
  assign _T_1030 = dut_io_coverage_115;
  assign _T_1031 = ~ dut_io_coverage_115;
  assign _T_1035 = {6'h0,SaturatingCounter_229_io_value};
  assign coverage_115 = {_T_1035,SaturatingCounter_230_io_value};
  assign _T_1037 = dut_io_coverage_116;
  assign _T_1038 = ~ dut_io_coverage_116;
  assign _T_1042 = {6'h0,SaturatingCounter_231_io_value};
  assign coverage_116 = {_T_1042,SaturatingCounter_232_io_value};
  assign _T_1044 = dut_io_coverage_117;
  assign _T_1045 = ~ dut_io_coverage_117;
  assign _T_1049 = {6'h0,SaturatingCounter_233_io_value};
  assign coverage_117 = {_T_1049,SaturatingCounter_234_io_value};
  assign _T_1051 = dut_io_coverage_118;
  assign _T_1052 = ~ dut_io_coverage_118;
  assign _T_1056 = {6'h0,SaturatingCounter_235_io_value};
  assign coverage_118 = {_T_1056,SaturatingCounter_236_io_value};
  assign _T_1058 = dut_io_coverage_119;
  assign _T_1059 = ~ dut_io_coverage_119;
  assign _T_1063 = {6'h0,SaturatingCounter_237_io_value};
  assign coverage_119 = {_T_1063,SaturatingCounter_238_io_value};
  assign _T_1065 = dut_io_coverage_120;
  assign _T_1066 = ~ dut_io_coverage_120;
  assign _T_1070 = {6'h0,SaturatingCounter_239_io_value};
  assign coverage_120 = {_T_1070,SaturatingCounter_240_io_value};
  assign _T_1072 = dut_io_coverage_121;
  assign _T_1073 = ~ dut_io_coverage_121;
  assign _T_1077 = {6'h0,SaturatingCounter_241_io_value};
  assign coverage_121 = {_T_1077,SaturatingCounter_242_io_value};
  assign _T_1079 = dut_io_coverage_122;
  assign _T_1080 = ~ dut_io_coverage_122;
  assign _T_1084 = {6'h0,SaturatingCounter_243_io_value};
  assign coverage_122 = {_T_1084,SaturatingCounter_244_io_value};
  assign _T_1086 = dut_io_coverage_123;
  assign _T_1087 = ~ dut_io_coverage_123;
  assign _T_1091 = {6'h0,SaturatingCounter_245_io_value};
  assign coverage_123 = {_T_1091,SaturatingCounter_246_io_value};
  assign _T_1093 = dut_io_coverage_124;
  assign _T_1094 = ~ dut_io_coverage_124;
  assign _T_1098 = {6'h0,SaturatingCounter_247_io_value};
  assign coverage_124 = {_T_1098,SaturatingCounter_248_io_value};
  assign _T_1100 = dut_io_coverage_125;
  assign _T_1101 = ~ dut_io_coverage_125;
  assign _T_1105 = {6'h0,SaturatingCounter_249_io_value};
  assign coverage_125 = {_T_1105,SaturatingCounter_250_io_value};
  assign _T_1107 = dut_io_coverage_126;
  assign _T_1108 = ~ dut_io_coverage_126;
  assign _T_1112 = {6'h0,SaturatingCounter_251_io_value};
  assign coverage_126 = {_T_1112,SaturatingCounter_252_io_value};
  assign _T_1114 = dut_io_coverage_127;
  assign _T_1115 = ~ dut_io_coverage_127;
  assign _T_1119 = {6'h0,SaturatingCounter_253_io_value};
  assign coverage_127 = {_T_1119,SaturatingCounter_254_io_value};
  assign _T_1121 = dut_io_coverage_128;
  assign _T_1122 = ~ dut_io_coverage_128;
  assign _T_1126 = {6'h0,SaturatingCounter_255_io_value};
  assign coverage_128 = {_T_1126,SaturatingCounter_256_io_value};
  assign _T_1128 = dut_io_coverage_129;
  assign _T_1129 = ~ dut_io_coverage_129;
  assign _T_1133 = {6'h0,SaturatingCounter_257_io_value};
  assign coverage_129 = {_T_1133,SaturatingCounter_258_io_value};
  assign _T_1135 = dut_io_coverage_130;
  assign _T_1136 = ~ dut_io_coverage_130;
  assign _T_1140 = {6'h0,SaturatingCounter_259_io_value};
  assign coverage_130 = {_T_1140,SaturatingCounter_260_io_value};
  assign _T_1142 = dut_io_coverage_131;
  assign _T_1143 = ~ dut_io_coverage_131;
  assign _T_1147 = {6'h0,SaturatingCounter_261_io_value};
  assign coverage_131 = {_T_1147,SaturatingCounter_262_io_value};
  assign _T_1149 = dut_io_coverage_132;
  assign _T_1150 = ~ dut_io_coverage_132;
  assign _T_1154 = {6'h0,SaturatingCounter_263_io_value};
  assign coverage_132 = {_T_1154,SaturatingCounter_264_io_value};
  assign _T_1156 = dut_io_coverage_133;
  assign _T_1157 = ~ dut_io_coverage_133;
  assign _T_1161 = {6'h0,SaturatingCounter_265_io_value};
  assign coverage_133 = {_T_1161,SaturatingCounter_266_io_value};
  assign _T_1163 = dut_io_coverage_134;
  assign _T_1164 = ~ dut_io_coverage_134;
  assign _T_1168 = {6'h0,SaturatingCounter_267_io_value};
  assign coverage_134 = {_T_1168,SaturatingCounter_268_io_value};
  assign _T_1170 = dut_io_coverage_135;
  assign _T_1171 = ~ dut_io_coverage_135;
  assign _T_1175 = {6'h0,SaturatingCounter_269_io_value};
  assign coverage_135 = {_T_1175,SaturatingCounter_270_io_value};
  assign _T_1177 = dut_io_coverage_136;
  assign _T_1178 = ~ dut_io_coverage_136;
  assign _T_1182 = {6'h0,SaturatingCounter_271_io_value};
  assign coverage_136 = {_T_1182,SaturatingCounter_272_io_value};
  assign _T_1184 = dut_io_coverage_137;
  assign _T_1185 = ~ dut_io_coverage_137;
  assign _T_1189 = {6'h0,SaturatingCounter_273_io_value};
  assign coverage_137 = {_T_1189,SaturatingCounter_274_io_value};
  assign _T_1191 = dut_io_coverage_138;
  assign _T_1192 = ~ dut_io_coverage_138;
  assign _T_1196 = {6'h0,SaturatingCounter_275_io_value};
  assign coverage_138 = {_T_1196,SaturatingCounter_276_io_value};
  assign _T_1198 = dut_io_coverage_139;
  assign _T_1199 = ~ dut_io_coverage_139;
  assign _T_1203 = {6'h0,SaturatingCounter_277_io_value};
  assign coverage_139 = {_T_1203,SaturatingCounter_278_io_value};
  assign _T_1205 = dut_io_coverage_140;
  assign _T_1206 = ~ dut_io_coverage_140;
  assign _T_1210 = {6'h0,SaturatingCounter_279_io_value};
  assign coverage_140 = {_T_1210,SaturatingCounter_280_io_value};
  assign _T_1212 = dut_io_coverage_141;
  assign _T_1213 = ~ dut_io_coverage_141;
  assign _T_1217 = {6'h0,SaturatingCounter_281_io_value};
  assign coverage_141 = {_T_1217,SaturatingCounter_282_io_value};
  assign _T_1219 = dut_io_coverage_142;
  assign _T_1220 = ~ dut_io_coverage_142;
  assign _T_1224 = {6'h0,SaturatingCounter_283_io_value};
  assign coverage_142 = {_T_1224,SaturatingCounter_284_io_value};
  assign _T_1226 = dut_io_coverage_143;
  assign _T_1227 = ~ dut_io_coverage_143;
  assign _T_1231 = {6'h0,SaturatingCounter_285_io_value};
  assign coverage_143 = {_T_1231,SaturatingCounter_286_io_value};
  assign _T_1233 = dut_io_coverage_144;
  assign _T_1234 = ~ dut_io_coverage_144;
  assign _T_1238 = {6'h0,SaturatingCounter_287_io_value};
  assign coverage_144 = {_T_1238,SaturatingCounter_288_io_value};
  assign _T_1240 = dut_io_coverage_145;
  assign _T_1241 = ~ dut_io_coverage_145;
  assign _T_1245 = {6'h0,SaturatingCounter_289_io_value};
  assign coverage_145 = {_T_1245,SaturatingCounter_290_io_value};
  assign _T_1247 = dut_io_coverage_146;
  assign _T_1248 = ~ dut_io_coverage_146;
  assign _T_1252 = {6'h0,SaturatingCounter_291_io_value};
  assign coverage_146 = {_T_1252,SaturatingCounter_292_io_value};
  assign _T_1254 = dut_io_coverage_147;
  assign _T_1255 = ~ dut_io_coverage_147;
  assign _T_1259 = {6'h0,SaturatingCounter_293_io_value};
  assign coverage_147 = {_T_1259,SaturatingCounter_294_io_value};
  assign _T_1261 = dut_io_coverage_148;
  assign _T_1262 = ~ dut_io_coverage_148;
  assign _T_1266 = {6'h0,SaturatingCounter_295_io_value};
  assign coverage_148 = {_T_1266,SaturatingCounter_296_io_value};
  assign _T_1268 = dut_io_coverage_149;
  assign _T_1269 = ~ dut_io_coverage_149;
  assign _T_1273 = {6'h0,SaturatingCounter_297_io_value};
  assign coverage_149 = {_T_1273,SaturatingCounter_298_io_value};
  assign _T_1275 = dut_io_coverage_150;
  assign _T_1276 = ~ dut_io_coverage_150;
  assign _T_1280 = {6'h0,SaturatingCounter_299_io_value};
  assign coverage_150 = {_T_1280,SaturatingCounter_300_io_value};
  assign _T_1282 = dut_io_coverage_151;
  assign _T_1283 = ~ dut_io_coverage_151;
  assign _T_1287 = {6'h0,SaturatingCounter_301_io_value};
  assign coverage_151 = {_T_1287,SaturatingCounter_302_io_value};
  assign _T_1289 = dut_io_coverage_152;
  assign _T_1290 = ~ dut_io_coverage_152;
  assign _T_1294 = {6'h0,SaturatingCounter_303_io_value};
  assign coverage_152 = {_T_1294,SaturatingCounter_304_io_value};
  assign _T_1296 = dut_io_coverage_153;
  assign _T_1297 = ~ dut_io_coverage_153;
  assign _T_1301 = {6'h0,SaturatingCounter_305_io_value};
  assign coverage_153 = {_T_1301,SaturatingCounter_306_io_value};
  assign _T_1303 = dut_io_coverage_154;
  assign _T_1304 = ~ dut_io_coverage_154;
  assign _T_1308 = {6'h0,SaturatingCounter_307_io_value};
  assign coverage_154 = {_T_1308,SaturatingCounter_308_io_value};
  assign _T_1310 = dut_io_coverage_155;
  assign _T_1311 = ~ dut_io_coverage_155;
  assign _T_1315 = {6'h0,SaturatingCounter_309_io_value};
  assign coverage_155 = {_T_1315,SaturatingCounter_310_io_value};
  assign _T_1317 = dut_io_coverage_156;
  assign _T_1318 = ~ dut_io_coverage_156;
  assign _T_1322 = {6'h0,SaturatingCounter_311_io_value};
  assign coverage_156 = {_T_1322,SaturatingCounter_312_io_value};
  assign _T_1324 = dut_io_coverage_157;
  assign _T_1325 = ~ dut_io_coverage_157;
  assign _T_1329 = {6'h0,SaturatingCounter_313_io_value};
  assign coverage_157 = {_T_1329,SaturatingCounter_314_io_value};
  assign _T_1331 = dut_io_coverage_158;
  assign _T_1332 = ~ dut_io_coverage_158;
  assign _T_1336 = {6'h0,SaturatingCounter_315_io_value};
  assign coverage_158 = {_T_1336,SaturatingCounter_316_io_value};
  assign _T_1338 = dut_io_coverage_159;
  assign _T_1339 = ~ dut_io_coverage_159;
  assign _T_1343 = {6'h0,SaturatingCounter_317_io_value};
  assign coverage_159 = {_T_1343,SaturatingCounter_318_io_value};
  assign _T_1345 = dut_io_coverage_160;
  assign _T_1346 = ~ dut_io_coverage_160;
  assign _T_1350 = {6'h0,SaturatingCounter_319_io_value};
  assign coverage_160 = {_T_1350,SaturatingCounter_320_io_value};
  assign _T_1352 = dut_io_coverage_161;
  assign _T_1353 = ~ dut_io_coverage_161;
  assign _T_1357 = {6'h0,SaturatingCounter_321_io_value};
  assign coverage_161 = {_T_1357,SaturatingCounter_322_io_value};
  assign _T_1359 = dut_io_coverage_162;
  assign _T_1360 = ~ dut_io_coverage_162;
  assign _T_1364 = {6'h0,SaturatingCounter_323_io_value};
  assign coverage_162 = {_T_1364,SaturatingCounter_324_io_value};
  assign _T_1366 = dut_io_coverage_163;
  assign _T_1367 = ~ dut_io_coverage_163;
  assign _T_1371 = {6'h0,SaturatingCounter_325_io_value};
  assign coverage_163 = {_T_1371,SaturatingCounter_326_io_value};
  assign _T_1373 = dut_io_coverage_164;
  assign _T_1374 = ~ dut_io_coverage_164;
  assign _T_1378 = {6'h0,SaturatingCounter_327_io_value};
  assign coverage_164 = {_T_1378,SaturatingCounter_328_io_value};
  assign _T_1380 = dut_io_coverage_165;
  assign _T_1381 = ~ dut_io_coverage_165;
  assign _T_1385 = {6'h0,SaturatingCounter_329_io_value};
  assign coverage_165 = {_T_1385,SaturatingCounter_330_io_value};
  assign _T_1387 = dut_io_coverage_166;
  assign _T_1388 = ~ dut_io_coverage_166;
  assign _T_1392 = {6'h0,SaturatingCounter_331_io_value};
  assign coverage_166 = {_T_1392,SaturatingCounter_332_io_value};
  assign _T_1394 = dut_io_coverage_167;
  assign _T_1395 = ~ dut_io_coverage_167;
  assign _T_1399 = {6'h0,SaturatingCounter_333_io_value};
  assign coverage_167 = {_T_1399,SaturatingCounter_334_io_value};
  assign _T_1401 = dut_io_coverage_168;
  assign _T_1402 = ~ dut_io_coverage_168;
  assign _T_1406 = {6'h0,SaturatingCounter_335_io_value};
  assign coverage_168 = {_T_1406,SaturatingCounter_336_io_value};
  assign _T_1408 = dut_io_coverage_169;
  assign _T_1409 = ~ dut_io_coverage_169;
  assign _T_1413 = {6'h0,SaturatingCounter_337_io_value};
  assign coverage_169 = {_T_1413,SaturatingCounter_338_io_value};
  assign _T_1415 = dut_io_coverage_170;
  assign _T_1416 = ~ dut_io_coverage_170;
  assign _T_1420 = {6'h0,SaturatingCounter_339_io_value};
  assign coverage_170 = {_T_1420,SaturatingCounter_340_io_value};
  assign _T_1422 = dut_io_coverage_171;
  assign _T_1423 = ~ dut_io_coverage_171;
  assign _T_1427 = {6'h0,SaturatingCounter_341_io_value};
  assign coverage_171 = {_T_1427,SaturatingCounter_342_io_value};
  assign _T_1429 = dut_io_coverage_172;
  assign _T_1430 = ~ dut_io_coverage_172;
  assign _T_1434 = {6'h0,SaturatingCounter_343_io_value};
  assign coverage_172 = {_T_1434,SaturatingCounter_344_io_value};
  assign _T_1436 = dut_io_coverage_173;
  assign _T_1437 = ~ dut_io_coverage_173;
  assign _T_1441 = {6'h0,SaturatingCounter_345_io_value};
  assign coverage_173 = {_T_1441,SaturatingCounter_346_io_value};
  assign _T_1443 = dut_io_coverage_174;
  assign _T_1444 = ~ dut_io_coverage_174;
  assign _T_1448 = {6'h0,SaturatingCounter_347_io_value};
  assign coverage_174 = {_T_1448,SaturatingCounter_348_io_value};
  assign _T_1450 = dut_io_coverage_175;
  assign _T_1451 = ~ dut_io_coverage_175;
  assign _T_1455 = {6'h0,SaturatingCounter_349_io_value};
  assign coverage_175 = {_T_1455,SaturatingCounter_350_io_value};
  assign _T_1457 = dut_io_coverage_176;
  assign _T_1458 = ~ dut_io_coverage_176;
  assign _T_1462 = {6'h0,SaturatingCounter_351_io_value};
  assign coverage_176 = {_T_1462,SaturatingCounter_352_io_value};
  assign _T_1464 = dut_io_coverage_177;
  assign _T_1465 = ~ dut_io_coverage_177;
  assign _T_1469 = {6'h0,SaturatingCounter_353_io_value};
  assign coverage_177 = {_T_1469,SaturatingCounter_354_io_value};
  assign _T_1471 = dut_io_coverage_178;
  assign _T_1472 = ~ dut_io_coverage_178;
  assign _T_1476 = {6'h0,SaturatingCounter_355_io_value};
  assign coverage_178 = {_T_1476,SaturatingCounter_356_io_value};
  assign _T_1478 = dut_io_coverage_179;
  assign _T_1479 = ~ dut_io_coverage_179;
  assign _T_1483 = {6'h0,SaturatingCounter_357_io_value};
  assign coverage_179 = {_T_1483,SaturatingCounter_358_io_value};
  assign _T_1485 = dut_io_coverage_180;
  assign _T_1486 = ~ dut_io_coverage_180;
  assign _T_1490 = {6'h0,SaturatingCounter_359_io_value};
  assign coverage_180 = {_T_1490,SaturatingCounter_360_io_value};
  assign _T_1492 = dut_io_coverage_181;
  assign _T_1493 = ~ dut_io_coverage_181;
  assign _T_1497 = {6'h0,SaturatingCounter_361_io_value};
  assign coverage_181 = {_T_1497,SaturatingCounter_362_io_value};
  assign _T_1499 = dut_io_coverage_182;
  assign _T_1500 = ~ dut_io_coverage_182;
  assign _T_1504 = {6'h0,SaturatingCounter_363_io_value};
  assign coverage_182 = {_T_1504,SaturatingCounter_364_io_value};
  assign _T_1506 = dut_io_coverage_183;
  assign _T_1507 = ~ dut_io_coverage_183;
  assign _T_1511 = {6'h0,SaturatingCounter_365_io_value};
  assign coverage_183 = {_T_1511,SaturatingCounter_366_io_value};
  assign _T_1513 = dut_io_coverage_184;
  assign _T_1514 = ~ dut_io_coverage_184;
  assign _T_1518 = {6'h0,SaturatingCounter_367_io_value};
  assign coverage_184 = {_T_1518,SaturatingCounter_368_io_value};
  assign _T_1520 = dut_io_coverage_185;
  assign _T_1521 = ~ dut_io_coverage_185;
  assign _T_1525 = {6'h0,SaturatingCounter_369_io_value};
  assign coverage_185 = {_T_1525,SaturatingCounter_370_io_value};
  assign _T_1527 = dut_io_coverage_186;
  assign _T_1528 = ~ dut_io_coverage_186;
  assign _T_1532 = {6'h0,SaturatingCounter_371_io_value};
  assign coverage_186 = {_T_1532,SaturatingCounter_372_io_value};
  assign _T_1534 = dut_io_coverage_187;
  assign _T_1535 = ~ dut_io_coverage_187;
  assign _T_1539 = {6'h0,SaturatingCounter_373_io_value};
  assign coverage_187 = {_T_1539,SaturatingCounter_374_io_value};
  assign _T_1541 = dut_io_coverage_188;
  assign _T_1542 = ~ dut_io_coverage_188;
  assign _T_1546 = {6'h0,SaturatingCounter_375_io_value};
  assign coverage_188 = {_T_1546,SaturatingCounter_376_io_value};
  assign _T_1548 = dut_io_coverage_189;
  assign _T_1549 = ~ dut_io_coverage_189;
  assign _T_1553 = {6'h0,SaturatingCounter_377_io_value};
  assign coverage_189 = {_T_1553,SaturatingCounter_378_io_value};
  assign _T_1555 = dut_io_coverage_190;
  assign _T_1556 = ~ dut_io_coverage_190;
  assign _T_1560 = {6'h0,SaturatingCounter_379_io_value};
  assign coverage_190 = {_T_1560,SaturatingCounter_380_io_value};
  assign _T_1562 = dut_io_coverage_191;
  assign _T_1563 = ~ dut_io_coverage_191;
  assign _T_1567 = {6'h0,SaturatingCounter_381_io_value};
  assign coverage_191 = {_T_1567,SaturatingCounter_382_io_value};
  assign io_coverage_bytes_0 = coverage_0;
  assign io_coverage_bytes_1 = coverage_1;
  assign io_coverage_bytes_2 = coverage_2;
  assign io_coverage_bytes_3 = coverage_3;
  assign io_coverage_bytes_4 = coverage_4;
  assign io_coverage_bytes_5 = coverage_5;
  assign io_coverage_bytes_6 = coverage_6;
  assign io_coverage_bytes_7 = coverage_7;
  assign io_coverage_bytes_8 = coverage_8;
  assign io_coverage_bytes_9 = coverage_9;
  assign io_coverage_bytes_10 = coverage_10;
  assign io_coverage_bytes_11 = coverage_11;
  assign io_coverage_bytes_12 = coverage_12;
  assign io_coverage_bytes_13 = coverage_13;
  assign io_coverage_bytes_14 = coverage_14;
  assign io_coverage_bytes_15 = coverage_15;
  assign io_coverage_bytes_16 = coverage_16;
  assign io_coverage_bytes_17 = coverage_17;
  assign io_coverage_bytes_18 = coverage_18;
  assign io_coverage_bytes_19 = coverage_19;
  assign io_coverage_bytes_20 = coverage_20;
  assign io_coverage_bytes_21 = coverage_21;
  assign io_coverage_bytes_22 = coverage_22;
  assign io_coverage_bytes_23 = coverage_23;
  assign io_coverage_bytes_24 = coverage_24;
  assign io_coverage_bytes_25 = coverage_25;
  assign io_coverage_bytes_26 = coverage_26;
  assign io_coverage_bytes_27 = coverage_27;
  assign io_coverage_bytes_28 = coverage_28;
  assign io_coverage_bytes_29 = coverage_29;
  assign io_coverage_bytes_30 = coverage_30;
  assign io_coverage_bytes_31 = coverage_31;
  assign io_coverage_bytes_32 = coverage_32;
  assign io_coverage_bytes_33 = coverage_33;
  assign io_coverage_bytes_34 = coverage_34;
  assign io_coverage_bytes_35 = coverage_35;
  assign io_coverage_bytes_36 = coverage_36;
  assign io_coverage_bytes_37 = coverage_37;
  assign io_coverage_bytes_38 = coverage_38;
  assign io_coverage_bytes_39 = coverage_39;
  assign io_coverage_bytes_40 = coverage_40;
  assign io_coverage_bytes_41 = coverage_41;
  assign io_coverage_bytes_42 = coverage_42;
  assign io_coverage_bytes_43 = coverage_43;
  assign io_coverage_bytes_44 = coverage_44;
  assign io_coverage_bytes_45 = coverage_45;
  assign io_coverage_bytes_46 = coverage_46;
  assign io_coverage_bytes_47 = coverage_47;
  assign io_coverage_bytes_48 = coverage_48;
  assign io_coverage_bytes_49 = coverage_49;
  assign io_coverage_bytes_50 = coverage_50;
  assign io_coverage_bytes_51 = coverage_51;
  assign io_coverage_bytes_52 = coverage_52;
  assign io_coverage_bytes_53 = coverage_53;
  assign io_coverage_bytes_54 = coverage_54;
  assign io_coverage_bytes_55 = coverage_55;
  assign io_coverage_bytes_56 = coverage_56;
  assign io_coverage_bytes_57 = coverage_57;
  assign io_coverage_bytes_58 = coverage_58;
  assign io_coverage_bytes_59 = coverage_59;
  assign io_coverage_bytes_60 = coverage_60;
  assign io_coverage_bytes_61 = coverage_61;
  assign io_coverage_bytes_62 = coverage_62;
  assign io_coverage_bytes_63 = coverage_63;
  assign io_coverage_bytes_64 = coverage_64;
  assign io_coverage_bytes_65 = coverage_65;
  assign io_coverage_bytes_66 = coverage_66;
  assign io_coverage_bytes_67 = coverage_67;
  assign io_coverage_bytes_68 = coverage_68;
  assign io_coverage_bytes_69 = coverage_69;
  assign io_coverage_bytes_70 = coverage_70;
  assign io_coverage_bytes_71 = coverage_71;
  assign io_coverage_bytes_72 = coverage_72;
  assign io_coverage_bytes_73 = coverage_73;
  assign io_coverage_bytes_74 = coverage_74;
  assign io_coverage_bytes_75 = coverage_75;
  assign io_coverage_bytes_76 = coverage_76;
  assign io_coverage_bytes_77 = coverage_77;
  assign io_coverage_bytes_78 = coverage_78;
  assign io_coverage_bytes_79 = coverage_79;
  assign io_coverage_bytes_80 = coverage_80;
  assign io_coverage_bytes_81 = coverage_81;
  assign io_coverage_bytes_82 = coverage_82;
  assign io_coverage_bytes_83 = coverage_83;
  assign io_coverage_bytes_84 = coverage_84;
  assign io_coverage_bytes_85 = coverage_85;
  assign io_coverage_bytes_86 = coverage_86;
  assign io_coverage_bytes_87 = coverage_87;
  assign io_coverage_bytes_88 = coverage_88;
  assign io_coverage_bytes_89 = coverage_89;
  assign io_coverage_bytes_90 = coverage_90;
  assign io_coverage_bytes_91 = coverage_91;
  assign io_coverage_bytes_92 = coverage_92;
  assign io_coverage_bytes_93 = coverage_93;
  assign io_coverage_bytes_94 = coverage_94;
  assign io_coverage_bytes_95 = coverage_95;
  assign io_coverage_bytes_96 = coverage_96;
  assign io_coverage_bytes_97 = coverage_97;
  assign io_coverage_bytes_98 = coverage_98;
  assign io_coverage_bytes_99 = coverage_99;
  assign io_coverage_bytes_100 = coverage_100;
  assign io_coverage_bytes_101 = coverage_101;
  assign io_coverage_bytes_102 = coverage_102;
  assign io_coverage_bytes_103 = coverage_103;
  assign io_coverage_bytes_104 = coverage_104;
  assign io_coverage_bytes_105 = coverage_105;
  assign io_coverage_bytes_106 = coverage_106;
  assign io_coverage_bytes_107 = coverage_107;
  assign io_coverage_bytes_108 = coverage_108;
  assign io_coverage_bytes_109 = coverage_109;
  assign io_coverage_bytes_110 = coverage_110;
  assign io_coverage_bytes_111 = coverage_111;
  assign io_coverage_bytes_112 = coverage_112;
  assign io_coverage_bytes_113 = coverage_113;
  assign io_coverage_bytes_114 = coverage_114;
  assign io_coverage_bytes_115 = coverage_115;
  assign io_coverage_bytes_116 = coverage_116;
  assign io_coverage_bytes_117 = coverage_117;
  assign io_coverage_bytes_118 = coverage_118;
  assign io_coverage_bytes_119 = coverage_119;
  assign io_coverage_bytes_120 = coverage_120;
  assign io_coverage_bytes_121 = coverage_121;
  assign io_coverage_bytes_122 = coverage_122;
  assign io_coverage_bytes_123 = coverage_123;
  assign io_coverage_bytes_124 = coverage_124;
  assign io_coverage_bytes_125 = coverage_125;
  assign io_coverage_bytes_126 = coverage_126;
  assign io_coverage_bytes_127 = coverage_127;
  assign io_coverage_bytes_128 = coverage_128;
  assign io_coverage_bytes_129 = coverage_129;
  assign io_coverage_bytes_130 = coverage_130;
  assign io_coverage_bytes_131 = coverage_131;
  assign io_coverage_bytes_132 = coverage_132;
  assign io_coverage_bytes_133 = coverage_133;
  assign io_coverage_bytes_134 = coverage_134;
  assign io_coverage_bytes_135 = coverage_135;
  assign io_coverage_bytes_136 = coverage_136;
  assign io_coverage_bytes_137 = coverage_137;
  assign io_coverage_bytes_138 = coverage_138;
  assign io_coverage_bytes_139 = coverage_139;
  assign io_coverage_bytes_140 = coverage_140;
  assign io_coverage_bytes_141 = coverage_141;
  assign io_coverage_bytes_142 = coverage_142;
  assign io_coverage_bytes_143 = coverage_143;
  assign io_coverage_bytes_144 = coverage_144;
  assign io_coverage_bytes_145 = coverage_145;
  assign io_coverage_bytes_146 = coverage_146;
  assign io_coverage_bytes_147 = coverage_147;
  assign io_coverage_bytes_148 = coverage_148;
  assign io_coverage_bytes_149 = coverage_149;
  assign io_coverage_bytes_150 = coverage_150;
  assign io_coverage_bytes_151 = coverage_151;
  assign io_coverage_bytes_152 = coverage_152;
  assign io_coverage_bytes_153 = coverage_153;
  assign io_coverage_bytes_154 = coverage_154;
  assign io_coverage_bytes_155 = coverage_155;
  assign io_coverage_bytes_156 = coverage_156;
  assign io_coverage_bytes_157 = coverage_157;
  assign io_coverage_bytes_158 = coverage_158;
  assign io_coverage_bytes_159 = coverage_159;
  assign io_coverage_bytes_160 = coverage_160;
  assign io_coverage_bytes_161 = coverage_161;
  assign io_coverage_bytes_162 = coverage_162;
  assign io_coverage_bytes_163 = coverage_163;
  assign io_coverage_bytes_164 = coverage_164;
  assign io_coverage_bytes_165 = coverage_165;
  assign io_coverage_bytes_166 = coverage_166;
  assign io_coverage_bytes_167 = coverage_167;
  assign io_coverage_bytes_168 = coverage_168;
  assign io_coverage_bytes_169 = coverage_169;
  assign io_coverage_bytes_170 = coverage_170;
  assign io_coverage_bytes_171 = coverage_171;
  assign io_coverage_bytes_172 = coverage_172;
  assign io_coverage_bytes_173 = coverage_173;
  assign io_coverage_bytes_174 = coverage_174;
  assign io_coverage_bytes_175 = coverage_175;
  assign io_coverage_bytes_176 = coverage_176;
  assign io_coverage_bytes_177 = coverage_177;
  assign io_coverage_bytes_178 = coverage_178;
  assign io_coverage_bytes_179 = coverage_179;
  assign io_coverage_bytes_180 = coverage_180;
  assign io_coverage_bytes_181 = coverage_181;
  assign io_coverage_bytes_182 = coverage_182;
  assign io_coverage_bytes_183 = coverage_183;
  assign io_coverage_bytes_184 = coverage_184;
  assign io_coverage_bytes_185 = coverage_185;
  assign io_coverage_bytes_186 = coverage_186;
  assign io_coverage_bytes_187 = coverage_187;
  assign io_coverage_bytes_188 = coverage_188;
  assign io_coverage_bytes_189 = coverage_189;
  assign io_coverage_bytes_190 = coverage_190;
  assign io_coverage_bytes_191 = coverage_191;
  assign io_coverage_bytes_192 = 8'h0;
  assign io_coverage_bytes_193 = 8'h0;
  assign io_coverage_bytes_194 = 8'h0;
  assign io_coverage_bytes_195 = 8'h0;
  assign io_coverage_bytes_196 = 8'h0;
  assign io_coverage_bytes_197 = 8'h0;
  assign dut_clock = clock;
  assign dut_reset = reset;
  assign dut_io_meta_reset = io_meta_reset;
  assign dut_io_inputs = _T_225;
  assign SaturatingCounter_clock = clock;
  assign SaturatingCounter_reset = reset;
  assign SaturatingCounter_io_enable = _T_227;
  assign SaturatingCounter_1_clock = clock;
  assign SaturatingCounter_1_reset = reset;
  assign SaturatingCounter_1_io_enable = _T_232;
  assign SaturatingCounter_2_clock = clock;
  assign SaturatingCounter_2_reset = reset;
  assign SaturatingCounter_2_io_enable = _T_233;
  assign SaturatingCounter_3_clock = clock;
  assign SaturatingCounter_3_reset = reset;
  assign SaturatingCounter_3_io_enable = _T_239;
  assign SaturatingCounter_4_clock = clock;
  assign SaturatingCounter_4_reset = reset;
  assign SaturatingCounter_4_io_enable = _T_240;
  assign SaturatingCounter_5_clock = clock;
  assign SaturatingCounter_5_reset = reset;
  assign SaturatingCounter_5_io_enable = _T_246;
  assign SaturatingCounter_6_clock = clock;
  assign SaturatingCounter_6_reset = reset;
  assign SaturatingCounter_6_io_enable = _T_247;
  assign SaturatingCounter_7_clock = clock;
  assign SaturatingCounter_7_reset = reset;
  assign SaturatingCounter_7_io_enable = _T_253;
  assign SaturatingCounter_8_clock = clock;
  assign SaturatingCounter_8_reset = reset;
  assign SaturatingCounter_8_io_enable = _T_254;
  assign SaturatingCounter_9_clock = clock;
  assign SaturatingCounter_9_reset = reset;
  assign SaturatingCounter_9_io_enable = _T_260;
  assign SaturatingCounter_10_clock = clock;
  assign SaturatingCounter_10_reset = reset;
  assign SaturatingCounter_10_io_enable = _T_261;
  assign SaturatingCounter_11_clock = clock;
  assign SaturatingCounter_11_reset = reset;
  assign SaturatingCounter_11_io_enable = _T_267;
  assign SaturatingCounter_12_clock = clock;
  assign SaturatingCounter_12_reset = reset;
  assign SaturatingCounter_12_io_enable = _T_268;
  assign SaturatingCounter_13_clock = clock;
  assign SaturatingCounter_13_reset = reset;
  assign SaturatingCounter_13_io_enable = _T_274;
  assign SaturatingCounter_14_clock = clock;
  assign SaturatingCounter_14_reset = reset;
  assign SaturatingCounter_14_io_enable = _T_275;
  assign SaturatingCounter_15_clock = clock;
  assign SaturatingCounter_15_reset = reset;
  assign SaturatingCounter_15_io_enable = _T_281;
  assign SaturatingCounter_16_clock = clock;
  assign SaturatingCounter_16_reset = reset;
  assign SaturatingCounter_16_io_enable = _T_282;
  assign SaturatingCounter_17_clock = clock;
  assign SaturatingCounter_17_reset = reset;
  assign SaturatingCounter_17_io_enable = _T_288;
  assign SaturatingCounter_18_clock = clock;
  assign SaturatingCounter_18_reset = reset;
  assign SaturatingCounter_18_io_enable = _T_289;
  assign SaturatingCounter_19_clock = clock;
  assign SaturatingCounter_19_reset = reset;
  assign SaturatingCounter_19_io_enable = _T_295;
  assign SaturatingCounter_20_clock = clock;
  assign SaturatingCounter_20_reset = reset;
  assign SaturatingCounter_20_io_enable = _T_296;
  assign SaturatingCounter_21_clock = clock;
  assign SaturatingCounter_21_reset = reset;
  assign SaturatingCounter_21_io_enable = _T_302;
  assign SaturatingCounter_22_clock = clock;
  assign SaturatingCounter_22_reset = reset;
  assign SaturatingCounter_22_io_enable = _T_303;
  assign SaturatingCounter_23_clock = clock;
  assign SaturatingCounter_23_reset = reset;
  assign SaturatingCounter_23_io_enable = _T_309;
  assign SaturatingCounter_24_clock = clock;
  assign SaturatingCounter_24_reset = reset;
  assign SaturatingCounter_24_io_enable = _T_310;
  assign SaturatingCounter_25_clock = clock;
  assign SaturatingCounter_25_reset = reset;
  assign SaturatingCounter_25_io_enable = _T_316;
  assign SaturatingCounter_26_clock = clock;
  assign SaturatingCounter_26_reset = reset;
  assign SaturatingCounter_26_io_enable = _T_317;
  assign SaturatingCounter_27_clock = clock;
  assign SaturatingCounter_27_reset = reset;
  assign SaturatingCounter_27_io_enable = _T_323;
  assign SaturatingCounter_28_clock = clock;
  assign SaturatingCounter_28_reset = reset;
  assign SaturatingCounter_28_io_enable = _T_324;
  assign SaturatingCounter_29_clock = clock;
  assign SaturatingCounter_29_reset = reset;
  assign SaturatingCounter_29_io_enable = _T_330;
  assign SaturatingCounter_30_clock = clock;
  assign SaturatingCounter_30_reset = reset;
  assign SaturatingCounter_30_io_enable = _T_331;
  assign SaturatingCounter_31_clock = clock;
  assign SaturatingCounter_31_reset = reset;
  assign SaturatingCounter_31_io_enable = _T_337;
  assign SaturatingCounter_32_clock = clock;
  assign SaturatingCounter_32_reset = reset;
  assign SaturatingCounter_32_io_enable = _T_338;
  assign SaturatingCounter_33_clock = clock;
  assign SaturatingCounter_33_reset = reset;
  assign SaturatingCounter_33_io_enable = _T_344;
  assign SaturatingCounter_34_clock = clock;
  assign SaturatingCounter_34_reset = reset;
  assign SaturatingCounter_34_io_enable = _T_345;
  assign SaturatingCounter_35_clock = clock;
  assign SaturatingCounter_35_reset = reset;
  assign SaturatingCounter_35_io_enable = _T_351;
  assign SaturatingCounter_36_clock = clock;
  assign SaturatingCounter_36_reset = reset;
  assign SaturatingCounter_36_io_enable = _T_352;
  assign SaturatingCounter_37_clock = clock;
  assign SaturatingCounter_37_reset = reset;
  assign SaturatingCounter_37_io_enable = _T_358;
  assign SaturatingCounter_38_clock = clock;
  assign SaturatingCounter_38_reset = reset;
  assign SaturatingCounter_38_io_enable = _T_359;
  assign SaturatingCounter_39_clock = clock;
  assign SaturatingCounter_39_reset = reset;
  assign SaturatingCounter_39_io_enable = _T_365;
  assign SaturatingCounter_40_clock = clock;
  assign SaturatingCounter_40_reset = reset;
  assign SaturatingCounter_40_io_enable = _T_366;
  assign SaturatingCounter_41_clock = clock;
  assign SaturatingCounter_41_reset = reset;
  assign SaturatingCounter_41_io_enable = _T_372;
  assign SaturatingCounter_42_clock = clock;
  assign SaturatingCounter_42_reset = reset;
  assign SaturatingCounter_42_io_enable = _T_373;
  assign SaturatingCounter_43_clock = clock;
  assign SaturatingCounter_43_reset = reset;
  assign SaturatingCounter_43_io_enable = _T_379;
  assign SaturatingCounter_44_clock = clock;
  assign SaturatingCounter_44_reset = reset;
  assign SaturatingCounter_44_io_enable = _T_380;
  assign SaturatingCounter_45_clock = clock;
  assign SaturatingCounter_45_reset = reset;
  assign SaturatingCounter_45_io_enable = _T_386;
  assign SaturatingCounter_46_clock = clock;
  assign SaturatingCounter_46_reset = reset;
  assign SaturatingCounter_46_io_enable = _T_387;
  assign SaturatingCounter_47_clock = clock;
  assign SaturatingCounter_47_reset = reset;
  assign SaturatingCounter_47_io_enable = _T_393;
  assign SaturatingCounter_48_clock = clock;
  assign SaturatingCounter_48_reset = reset;
  assign SaturatingCounter_48_io_enable = _T_394;
  assign SaturatingCounter_49_clock = clock;
  assign SaturatingCounter_49_reset = reset;
  assign SaturatingCounter_49_io_enable = _T_400;
  assign SaturatingCounter_50_clock = clock;
  assign SaturatingCounter_50_reset = reset;
  assign SaturatingCounter_50_io_enable = _T_401;
  assign SaturatingCounter_51_clock = clock;
  assign SaturatingCounter_51_reset = reset;
  assign SaturatingCounter_51_io_enable = _T_407;
  assign SaturatingCounter_52_clock = clock;
  assign SaturatingCounter_52_reset = reset;
  assign SaturatingCounter_52_io_enable = _T_408;
  assign SaturatingCounter_53_clock = clock;
  assign SaturatingCounter_53_reset = reset;
  assign SaturatingCounter_53_io_enable = _T_414;
  assign SaturatingCounter_54_clock = clock;
  assign SaturatingCounter_54_reset = reset;
  assign SaturatingCounter_54_io_enable = _T_415;
  assign SaturatingCounter_55_clock = clock;
  assign SaturatingCounter_55_reset = reset;
  assign SaturatingCounter_55_io_enable = _T_421;
  assign SaturatingCounter_56_clock = clock;
  assign SaturatingCounter_56_reset = reset;
  assign SaturatingCounter_56_io_enable = _T_422;
  assign SaturatingCounter_57_clock = clock;
  assign SaturatingCounter_57_reset = reset;
  assign SaturatingCounter_57_io_enable = _T_428;
  assign SaturatingCounter_58_clock = clock;
  assign SaturatingCounter_58_reset = reset;
  assign SaturatingCounter_58_io_enable = _T_429;
  assign SaturatingCounter_59_clock = clock;
  assign SaturatingCounter_59_reset = reset;
  assign SaturatingCounter_59_io_enable = _T_435;
  assign SaturatingCounter_60_clock = clock;
  assign SaturatingCounter_60_reset = reset;
  assign SaturatingCounter_60_io_enable = _T_436;
  assign SaturatingCounter_61_clock = clock;
  assign SaturatingCounter_61_reset = reset;
  assign SaturatingCounter_61_io_enable = _T_442;
  assign SaturatingCounter_62_clock = clock;
  assign SaturatingCounter_62_reset = reset;
  assign SaturatingCounter_62_io_enable = _T_443;
  assign SaturatingCounter_63_clock = clock;
  assign SaturatingCounter_63_reset = reset;
  assign SaturatingCounter_63_io_enable = _T_449;
  assign SaturatingCounter_64_clock = clock;
  assign SaturatingCounter_64_reset = reset;
  assign SaturatingCounter_64_io_enable = _T_450;
  assign SaturatingCounter_65_clock = clock;
  assign SaturatingCounter_65_reset = reset;
  assign SaturatingCounter_65_io_enable = _T_456;
  assign SaturatingCounter_66_clock = clock;
  assign SaturatingCounter_66_reset = reset;
  assign SaturatingCounter_66_io_enable = _T_457;
  assign SaturatingCounter_67_clock = clock;
  assign SaturatingCounter_67_reset = reset;
  assign SaturatingCounter_67_io_enable = _T_463;
  assign SaturatingCounter_68_clock = clock;
  assign SaturatingCounter_68_reset = reset;
  assign SaturatingCounter_68_io_enable = _T_464;
  assign SaturatingCounter_69_clock = clock;
  assign SaturatingCounter_69_reset = reset;
  assign SaturatingCounter_69_io_enable = _T_470;
  assign SaturatingCounter_70_clock = clock;
  assign SaturatingCounter_70_reset = reset;
  assign SaturatingCounter_70_io_enable = _T_471;
  assign SaturatingCounter_71_clock = clock;
  assign SaturatingCounter_71_reset = reset;
  assign SaturatingCounter_71_io_enable = _T_477;
  assign SaturatingCounter_72_clock = clock;
  assign SaturatingCounter_72_reset = reset;
  assign SaturatingCounter_72_io_enable = _T_478;
  assign SaturatingCounter_73_clock = clock;
  assign SaturatingCounter_73_reset = reset;
  assign SaturatingCounter_73_io_enable = _T_484;
  assign SaturatingCounter_74_clock = clock;
  assign SaturatingCounter_74_reset = reset;
  assign SaturatingCounter_74_io_enable = _T_485;
  assign SaturatingCounter_75_clock = clock;
  assign SaturatingCounter_75_reset = reset;
  assign SaturatingCounter_75_io_enable = _T_491;
  assign SaturatingCounter_76_clock = clock;
  assign SaturatingCounter_76_reset = reset;
  assign SaturatingCounter_76_io_enable = _T_492;
  assign SaturatingCounter_77_clock = clock;
  assign SaturatingCounter_77_reset = reset;
  assign SaturatingCounter_77_io_enable = _T_498;
  assign SaturatingCounter_78_clock = clock;
  assign SaturatingCounter_78_reset = reset;
  assign SaturatingCounter_78_io_enable = _T_499;
  assign SaturatingCounter_79_clock = clock;
  assign SaturatingCounter_79_reset = reset;
  assign SaturatingCounter_79_io_enable = _T_505;
  assign SaturatingCounter_80_clock = clock;
  assign SaturatingCounter_80_reset = reset;
  assign SaturatingCounter_80_io_enable = _T_506;
  assign SaturatingCounter_81_clock = clock;
  assign SaturatingCounter_81_reset = reset;
  assign SaturatingCounter_81_io_enable = _T_512;
  assign SaturatingCounter_82_clock = clock;
  assign SaturatingCounter_82_reset = reset;
  assign SaturatingCounter_82_io_enable = _T_513;
  assign SaturatingCounter_83_clock = clock;
  assign SaturatingCounter_83_reset = reset;
  assign SaturatingCounter_83_io_enable = _T_519;
  assign SaturatingCounter_84_clock = clock;
  assign SaturatingCounter_84_reset = reset;
  assign SaturatingCounter_84_io_enable = _T_520;
  assign SaturatingCounter_85_clock = clock;
  assign SaturatingCounter_85_reset = reset;
  assign SaturatingCounter_85_io_enable = _T_526;
  assign SaturatingCounter_86_clock = clock;
  assign SaturatingCounter_86_reset = reset;
  assign SaturatingCounter_86_io_enable = _T_527;
  assign SaturatingCounter_87_clock = clock;
  assign SaturatingCounter_87_reset = reset;
  assign SaturatingCounter_87_io_enable = _T_533;
  assign SaturatingCounter_88_clock = clock;
  assign SaturatingCounter_88_reset = reset;
  assign SaturatingCounter_88_io_enable = _T_534;
  assign SaturatingCounter_89_clock = clock;
  assign SaturatingCounter_89_reset = reset;
  assign SaturatingCounter_89_io_enable = _T_540;
  assign SaturatingCounter_90_clock = clock;
  assign SaturatingCounter_90_reset = reset;
  assign SaturatingCounter_90_io_enable = _T_541;
  assign SaturatingCounter_91_clock = clock;
  assign SaturatingCounter_91_reset = reset;
  assign SaturatingCounter_91_io_enable = _T_547;
  assign SaturatingCounter_92_clock = clock;
  assign SaturatingCounter_92_reset = reset;
  assign SaturatingCounter_92_io_enable = _T_548;
  assign SaturatingCounter_93_clock = clock;
  assign SaturatingCounter_93_reset = reset;
  assign SaturatingCounter_93_io_enable = _T_554;
  assign SaturatingCounter_94_clock = clock;
  assign SaturatingCounter_94_reset = reset;
  assign SaturatingCounter_94_io_enable = _T_555;
  assign SaturatingCounter_95_clock = clock;
  assign SaturatingCounter_95_reset = reset;
  assign SaturatingCounter_95_io_enable = _T_561;
  assign SaturatingCounter_96_clock = clock;
  assign SaturatingCounter_96_reset = reset;
  assign SaturatingCounter_96_io_enable = _T_562;
  assign SaturatingCounter_97_clock = clock;
  assign SaturatingCounter_97_reset = reset;
  assign SaturatingCounter_97_io_enable = _T_568;
  assign SaturatingCounter_98_clock = clock;
  assign SaturatingCounter_98_reset = reset;
  assign SaturatingCounter_98_io_enable = _T_569;
  assign SaturatingCounter_99_clock = clock;
  assign SaturatingCounter_99_reset = reset;
  assign SaturatingCounter_99_io_enable = _T_575;
  assign SaturatingCounter_100_clock = clock;
  assign SaturatingCounter_100_reset = reset;
  assign SaturatingCounter_100_io_enable = _T_576;
  assign SaturatingCounter_101_clock = clock;
  assign SaturatingCounter_101_reset = reset;
  assign SaturatingCounter_101_io_enable = _T_582;
  assign SaturatingCounter_102_clock = clock;
  assign SaturatingCounter_102_reset = reset;
  assign SaturatingCounter_102_io_enable = _T_583;
  assign SaturatingCounter_103_clock = clock;
  assign SaturatingCounter_103_reset = reset;
  assign SaturatingCounter_103_io_enable = _T_589;
  assign SaturatingCounter_104_clock = clock;
  assign SaturatingCounter_104_reset = reset;
  assign SaturatingCounter_104_io_enable = _T_590;
  assign SaturatingCounter_105_clock = clock;
  assign SaturatingCounter_105_reset = reset;
  assign SaturatingCounter_105_io_enable = _T_596;
  assign SaturatingCounter_106_clock = clock;
  assign SaturatingCounter_106_reset = reset;
  assign SaturatingCounter_106_io_enable = _T_597;
  assign SaturatingCounter_107_clock = clock;
  assign SaturatingCounter_107_reset = reset;
  assign SaturatingCounter_107_io_enable = _T_603;
  assign SaturatingCounter_108_clock = clock;
  assign SaturatingCounter_108_reset = reset;
  assign SaturatingCounter_108_io_enable = _T_604;
  assign SaturatingCounter_109_clock = clock;
  assign SaturatingCounter_109_reset = reset;
  assign SaturatingCounter_109_io_enable = _T_610;
  assign SaturatingCounter_110_clock = clock;
  assign SaturatingCounter_110_reset = reset;
  assign SaturatingCounter_110_io_enable = _T_611;
  assign SaturatingCounter_111_clock = clock;
  assign SaturatingCounter_111_reset = reset;
  assign SaturatingCounter_111_io_enable = _T_617;
  assign SaturatingCounter_112_clock = clock;
  assign SaturatingCounter_112_reset = reset;
  assign SaturatingCounter_112_io_enable = _T_618;
  assign SaturatingCounter_113_clock = clock;
  assign SaturatingCounter_113_reset = reset;
  assign SaturatingCounter_113_io_enable = _T_624;
  assign SaturatingCounter_114_clock = clock;
  assign SaturatingCounter_114_reset = reset;
  assign SaturatingCounter_114_io_enable = _T_625;
  assign SaturatingCounter_115_clock = clock;
  assign SaturatingCounter_115_reset = reset;
  assign SaturatingCounter_115_io_enable = _T_631;
  assign SaturatingCounter_116_clock = clock;
  assign SaturatingCounter_116_reset = reset;
  assign SaturatingCounter_116_io_enable = _T_632;
  assign SaturatingCounter_117_clock = clock;
  assign SaturatingCounter_117_reset = reset;
  assign SaturatingCounter_117_io_enable = _T_638;
  assign SaturatingCounter_118_clock = clock;
  assign SaturatingCounter_118_reset = reset;
  assign SaturatingCounter_118_io_enable = _T_639;
  assign SaturatingCounter_119_clock = clock;
  assign SaturatingCounter_119_reset = reset;
  assign SaturatingCounter_119_io_enable = _T_645;
  assign SaturatingCounter_120_clock = clock;
  assign SaturatingCounter_120_reset = reset;
  assign SaturatingCounter_120_io_enable = _T_646;
  assign SaturatingCounter_121_clock = clock;
  assign SaturatingCounter_121_reset = reset;
  assign SaturatingCounter_121_io_enable = _T_652;
  assign SaturatingCounter_122_clock = clock;
  assign SaturatingCounter_122_reset = reset;
  assign SaturatingCounter_122_io_enable = _T_653;
  assign SaturatingCounter_123_clock = clock;
  assign SaturatingCounter_123_reset = reset;
  assign SaturatingCounter_123_io_enable = _T_659;
  assign SaturatingCounter_124_clock = clock;
  assign SaturatingCounter_124_reset = reset;
  assign SaturatingCounter_124_io_enable = _T_660;
  assign SaturatingCounter_125_clock = clock;
  assign SaturatingCounter_125_reset = reset;
  assign SaturatingCounter_125_io_enable = _T_666;
  assign SaturatingCounter_126_clock = clock;
  assign SaturatingCounter_126_reset = reset;
  assign SaturatingCounter_126_io_enable = _T_667;
  assign SaturatingCounter_127_clock = clock;
  assign SaturatingCounter_127_reset = reset;
  assign SaturatingCounter_127_io_enable = _T_673;
  assign SaturatingCounter_128_clock = clock;
  assign SaturatingCounter_128_reset = reset;
  assign SaturatingCounter_128_io_enable = _T_674;
  assign SaturatingCounter_129_clock = clock;
  assign SaturatingCounter_129_reset = reset;
  assign SaturatingCounter_129_io_enable = _T_680;
  assign SaturatingCounter_130_clock = clock;
  assign SaturatingCounter_130_reset = reset;
  assign SaturatingCounter_130_io_enable = _T_681;
  assign SaturatingCounter_131_clock = clock;
  assign SaturatingCounter_131_reset = reset;
  assign SaturatingCounter_131_io_enable = _T_687;
  assign SaturatingCounter_132_clock = clock;
  assign SaturatingCounter_132_reset = reset;
  assign SaturatingCounter_132_io_enable = _T_688;
  assign SaturatingCounter_133_clock = clock;
  assign SaturatingCounter_133_reset = reset;
  assign SaturatingCounter_133_io_enable = _T_694;
  assign SaturatingCounter_134_clock = clock;
  assign SaturatingCounter_134_reset = reset;
  assign SaturatingCounter_134_io_enable = _T_695;
  assign SaturatingCounter_135_clock = clock;
  assign SaturatingCounter_135_reset = reset;
  assign SaturatingCounter_135_io_enable = _T_701;
  assign SaturatingCounter_136_clock = clock;
  assign SaturatingCounter_136_reset = reset;
  assign SaturatingCounter_136_io_enable = _T_702;
  assign SaturatingCounter_137_clock = clock;
  assign SaturatingCounter_137_reset = reset;
  assign SaturatingCounter_137_io_enable = _T_708;
  assign SaturatingCounter_138_clock = clock;
  assign SaturatingCounter_138_reset = reset;
  assign SaturatingCounter_138_io_enable = _T_709;
  assign SaturatingCounter_139_clock = clock;
  assign SaturatingCounter_139_reset = reset;
  assign SaturatingCounter_139_io_enable = _T_715;
  assign SaturatingCounter_140_clock = clock;
  assign SaturatingCounter_140_reset = reset;
  assign SaturatingCounter_140_io_enable = _T_716;
  assign SaturatingCounter_141_clock = clock;
  assign SaturatingCounter_141_reset = reset;
  assign SaturatingCounter_141_io_enable = _T_722;
  assign SaturatingCounter_142_clock = clock;
  assign SaturatingCounter_142_reset = reset;
  assign SaturatingCounter_142_io_enable = _T_723;
  assign SaturatingCounter_143_clock = clock;
  assign SaturatingCounter_143_reset = reset;
  assign SaturatingCounter_143_io_enable = _T_729;
  assign SaturatingCounter_144_clock = clock;
  assign SaturatingCounter_144_reset = reset;
  assign SaturatingCounter_144_io_enable = _T_730;
  assign SaturatingCounter_145_clock = clock;
  assign SaturatingCounter_145_reset = reset;
  assign SaturatingCounter_145_io_enable = _T_736;
  assign SaturatingCounter_146_clock = clock;
  assign SaturatingCounter_146_reset = reset;
  assign SaturatingCounter_146_io_enable = _T_737;
  assign SaturatingCounter_147_clock = clock;
  assign SaturatingCounter_147_reset = reset;
  assign SaturatingCounter_147_io_enable = _T_743;
  assign SaturatingCounter_148_clock = clock;
  assign SaturatingCounter_148_reset = reset;
  assign SaturatingCounter_148_io_enable = _T_744;
  assign SaturatingCounter_149_clock = clock;
  assign SaturatingCounter_149_reset = reset;
  assign SaturatingCounter_149_io_enable = _T_750;
  assign SaturatingCounter_150_clock = clock;
  assign SaturatingCounter_150_reset = reset;
  assign SaturatingCounter_150_io_enable = _T_751;
  assign SaturatingCounter_151_clock = clock;
  assign SaturatingCounter_151_reset = reset;
  assign SaturatingCounter_151_io_enable = _T_757;
  assign SaturatingCounter_152_clock = clock;
  assign SaturatingCounter_152_reset = reset;
  assign SaturatingCounter_152_io_enable = _T_758;
  assign SaturatingCounter_153_clock = clock;
  assign SaturatingCounter_153_reset = reset;
  assign SaturatingCounter_153_io_enable = _T_764;
  assign SaturatingCounter_154_clock = clock;
  assign SaturatingCounter_154_reset = reset;
  assign SaturatingCounter_154_io_enable = _T_765;
  assign SaturatingCounter_155_clock = clock;
  assign SaturatingCounter_155_reset = reset;
  assign SaturatingCounter_155_io_enable = _T_771;
  assign SaturatingCounter_156_clock = clock;
  assign SaturatingCounter_156_reset = reset;
  assign SaturatingCounter_156_io_enable = _T_772;
  assign SaturatingCounter_157_clock = clock;
  assign SaturatingCounter_157_reset = reset;
  assign SaturatingCounter_157_io_enable = _T_778;
  assign SaturatingCounter_158_clock = clock;
  assign SaturatingCounter_158_reset = reset;
  assign SaturatingCounter_158_io_enable = _T_779;
  assign SaturatingCounter_159_clock = clock;
  assign SaturatingCounter_159_reset = reset;
  assign SaturatingCounter_159_io_enable = _T_785;
  assign SaturatingCounter_160_clock = clock;
  assign SaturatingCounter_160_reset = reset;
  assign SaturatingCounter_160_io_enable = _T_786;
  assign SaturatingCounter_161_clock = clock;
  assign SaturatingCounter_161_reset = reset;
  assign SaturatingCounter_161_io_enable = _T_792;
  assign SaturatingCounter_162_clock = clock;
  assign SaturatingCounter_162_reset = reset;
  assign SaturatingCounter_162_io_enable = _T_793;
  assign SaturatingCounter_163_clock = clock;
  assign SaturatingCounter_163_reset = reset;
  assign SaturatingCounter_163_io_enable = _T_799;
  assign SaturatingCounter_164_clock = clock;
  assign SaturatingCounter_164_reset = reset;
  assign SaturatingCounter_164_io_enable = _T_800;
  assign SaturatingCounter_165_clock = clock;
  assign SaturatingCounter_165_reset = reset;
  assign SaturatingCounter_165_io_enable = _T_806;
  assign SaturatingCounter_166_clock = clock;
  assign SaturatingCounter_166_reset = reset;
  assign SaturatingCounter_166_io_enable = _T_807;
  assign SaturatingCounter_167_clock = clock;
  assign SaturatingCounter_167_reset = reset;
  assign SaturatingCounter_167_io_enable = _T_813;
  assign SaturatingCounter_168_clock = clock;
  assign SaturatingCounter_168_reset = reset;
  assign SaturatingCounter_168_io_enable = _T_814;
  assign SaturatingCounter_169_clock = clock;
  assign SaturatingCounter_169_reset = reset;
  assign SaturatingCounter_169_io_enable = _T_820;
  assign SaturatingCounter_170_clock = clock;
  assign SaturatingCounter_170_reset = reset;
  assign SaturatingCounter_170_io_enable = _T_821;
  assign SaturatingCounter_171_clock = clock;
  assign SaturatingCounter_171_reset = reset;
  assign SaturatingCounter_171_io_enable = _T_827;
  assign SaturatingCounter_172_clock = clock;
  assign SaturatingCounter_172_reset = reset;
  assign SaturatingCounter_172_io_enable = _T_828;
  assign SaturatingCounter_173_clock = clock;
  assign SaturatingCounter_173_reset = reset;
  assign SaturatingCounter_173_io_enable = _T_834;
  assign SaturatingCounter_174_clock = clock;
  assign SaturatingCounter_174_reset = reset;
  assign SaturatingCounter_174_io_enable = _T_835;
  assign SaturatingCounter_175_clock = clock;
  assign SaturatingCounter_175_reset = reset;
  assign SaturatingCounter_175_io_enable = _T_841;
  assign SaturatingCounter_176_clock = clock;
  assign SaturatingCounter_176_reset = reset;
  assign SaturatingCounter_176_io_enable = _T_842;
  assign SaturatingCounter_177_clock = clock;
  assign SaturatingCounter_177_reset = reset;
  assign SaturatingCounter_177_io_enable = _T_848;
  assign SaturatingCounter_178_clock = clock;
  assign SaturatingCounter_178_reset = reset;
  assign SaturatingCounter_178_io_enable = _T_849;
  assign SaturatingCounter_179_clock = clock;
  assign SaturatingCounter_179_reset = reset;
  assign SaturatingCounter_179_io_enable = _T_855;
  assign SaturatingCounter_180_clock = clock;
  assign SaturatingCounter_180_reset = reset;
  assign SaturatingCounter_180_io_enable = _T_856;
  assign SaturatingCounter_181_clock = clock;
  assign SaturatingCounter_181_reset = reset;
  assign SaturatingCounter_181_io_enable = _T_862;
  assign SaturatingCounter_182_clock = clock;
  assign SaturatingCounter_182_reset = reset;
  assign SaturatingCounter_182_io_enable = _T_863;
  assign SaturatingCounter_183_clock = clock;
  assign SaturatingCounter_183_reset = reset;
  assign SaturatingCounter_183_io_enable = _T_869;
  assign SaturatingCounter_184_clock = clock;
  assign SaturatingCounter_184_reset = reset;
  assign SaturatingCounter_184_io_enable = _T_870;
  assign SaturatingCounter_185_clock = clock;
  assign SaturatingCounter_185_reset = reset;
  assign SaturatingCounter_185_io_enable = _T_876;
  assign SaturatingCounter_186_clock = clock;
  assign SaturatingCounter_186_reset = reset;
  assign SaturatingCounter_186_io_enable = _T_877;
  assign SaturatingCounter_187_clock = clock;
  assign SaturatingCounter_187_reset = reset;
  assign SaturatingCounter_187_io_enable = _T_883;
  assign SaturatingCounter_188_clock = clock;
  assign SaturatingCounter_188_reset = reset;
  assign SaturatingCounter_188_io_enable = _T_884;
  assign SaturatingCounter_189_clock = clock;
  assign SaturatingCounter_189_reset = reset;
  assign SaturatingCounter_189_io_enable = _T_890;
  assign SaturatingCounter_190_clock = clock;
  assign SaturatingCounter_190_reset = reset;
  assign SaturatingCounter_190_io_enable = _T_891;
  assign SaturatingCounter_191_clock = clock;
  assign SaturatingCounter_191_reset = reset;
  assign SaturatingCounter_191_io_enable = _T_897;
  assign SaturatingCounter_192_clock = clock;
  assign SaturatingCounter_192_reset = reset;
  assign SaturatingCounter_192_io_enable = _T_898;
  assign SaturatingCounter_193_clock = clock;
  assign SaturatingCounter_193_reset = reset;
  assign SaturatingCounter_193_io_enable = _T_904;
  assign SaturatingCounter_194_clock = clock;
  assign SaturatingCounter_194_reset = reset;
  assign SaturatingCounter_194_io_enable = _T_905;
  assign SaturatingCounter_195_clock = clock;
  assign SaturatingCounter_195_reset = reset;
  assign SaturatingCounter_195_io_enable = _T_911;
  assign SaturatingCounter_196_clock = clock;
  assign SaturatingCounter_196_reset = reset;
  assign SaturatingCounter_196_io_enable = _T_912;
  assign SaturatingCounter_197_clock = clock;
  assign SaturatingCounter_197_reset = reset;
  assign SaturatingCounter_197_io_enable = _T_918;
  assign SaturatingCounter_198_clock = clock;
  assign SaturatingCounter_198_reset = reset;
  assign SaturatingCounter_198_io_enable = _T_919;
  assign SaturatingCounter_199_clock = clock;
  assign SaturatingCounter_199_reset = reset;
  assign SaturatingCounter_199_io_enable = _T_925;
  assign SaturatingCounter_200_clock = clock;
  assign SaturatingCounter_200_reset = reset;
  assign SaturatingCounter_200_io_enable = _T_926;
  assign SaturatingCounter_201_clock = clock;
  assign SaturatingCounter_201_reset = reset;
  assign SaturatingCounter_201_io_enable = _T_932;
  assign SaturatingCounter_202_clock = clock;
  assign SaturatingCounter_202_reset = reset;
  assign SaturatingCounter_202_io_enable = _T_933;
  assign SaturatingCounter_203_clock = clock;
  assign SaturatingCounter_203_reset = reset;
  assign SaturatingCounter_203_io_enable = _T_939;
  assign SaturatingCounter_204_clock = clock;
  assign SaturatingCounter_204_reset = reset;
  assign SaturatingCounter_204_io_enable = _T_940;
  assign SaturatingCounter_205_clock = clock;
  assign SaturatingCounter_205_reset = reset;
  assign SaturatingCounter_205_io_enable = _T_946;
  assign SaturatingCounter_206_clock = clock;
  assign SaturatingCounter_206_reset = reset;
  assign SaturatingCounter_206_io_enable = _T_947;
  assign SaturatingCounter_207_clock = clock;
  assign SaturatingCounter_207_reset = reset;
  assign SaturatingCounter_207_io_enable = _T_953;
  assign SaturatingCounter_208_clock = clock;
  assign SaturatingCounter_208_reset = reset;
  assign SaturatingCounter_208_io_enable = _T_954;
  assign SaturatingCounter_209_clock = clock;
  assign SaturatingCounter_209_reset = reset;
  assign SaturatingCounter_209_io_enable = _T_960;
  assign SaturatingCounter_210_clock = clock;
  assign SaturatingCounter_210_reset = reset;
  assign SaturatingCounter_210_io_enable = _T_961;
  assign SaturatingCounter_211_clock = clock;
  assign SaturatingCounter_211_reset = reset;
  assign SaturatingCounter_211_io_enable = _T_967;
  assign SaturatingCounter_212_clock = clock;
  assign SaturatingCounter_212_reset = reset;
  assign SaturatingCounter_212_io_enable = _T_968;
  assign SaturatingCounter_213_clock = clock;
  assign SaturatingCounter_213_reset = reset;
  assign SaturatingCounter_213_io_enable = _T_974;
  assign SaturatingCounter_214_clock = clock;
  assign SaturatingCounter_214_reset = reset;
  assign SaturatingCounter_214_io_enable = _T_975;
  assign SaturatingCounter_215_clock = clock;
  assign SaturatingCounter_215_reset = reset;
  assign SaturatingCounter_215_io_enable = _T_981;
  assign SaturatingCounter_216_clock = clock;
  assign SaturatingCounter_216_reset = reset;
  assign SaturatingCounter_216_io_enable = _T_982;
  assign SaturatingCounter_217_clock = clock;
  assign SaturatingCounter_217_reset = reset;
  assign SaturatingCounter_217_io_enable = _T_988;
  assign SaturatingCounter_218_clock = clock;
  assign SaturatingCounter_218_reset = reset;
  assign SaturatingCounter_218_io_enable = _T_989;
  assign SaturatingCounter_219_clock = clock;
  assign SaturatingCounter_219_reset = reset;
  assign SaturatingCounter_219_io_enable = _T_995;
  assign SaturatingCounter_220_clock = clock;
  assign SaturatingCounter_220_reset = reset;
  assign SaturatingCounter_220_io_enable = _T_996;
  assign SaturatingCounter_221_clock = clock;
  assign SaturatingCounter_221_reset = reset;
  assign SaturatingCounter_221_io_enable = _T_1002;
  assign SaturatingCounter_222_clock = clock;
  assign SaturatingCounter_222_reset = reset;
  assign SaturatingCounter_222_io_enable = _T_1003;
  assign SaturatingCounter_223_clock = clock;
  assign SaturatingCounter_223_reset = reset;
  assign SaturatingCounter_223_io_enable = _T_1009;
  assign SaturatingCounter_224_clock = clock;
  assign SaturatingCounter_224_reset = reset;
  assign SaturatingCounter_224_io_enable = _T_1010;
  assign SaturatingCounter_225_clock = clock;
  assign SaturatingCounter_225_reset = reset;
  assign SaturatingCounter_225_io_enable = _T_1016;
  assign SaturatingCounter_226_clock = clock;
  assign SaturatingCounter_226_reset = reset;
  assign SaturatingCounter_226_io_enable = _T_1017;
  assign SaturatingCounter_227_clock = clock;
  assign SaturatingCounter_227_reset = reset;
  assign SaturatingCounter_227_io_enable = _T_1023;
  assign SaturatingCounter_228_clock = clock;
  assign SaturatingCounter_228_reset = reset;
  assign SaturatingCounter_228_io_enable = _T_1024;
  assign SaturatingCounter_229_clock = clock;
  assign SaturatingCounter_229_reset = reset;
  assign SaturatingCounter_229_io_enable = _T_1030;
  assign SaturatingCounter_230_clock = clock;
  assign SaturatingCounter_230_reset = reset;
  assign SaturatingCounter_230_io_enable = _T_1031;
  assign SaturatingCounter_231_clock = clock;
  assign SaturatingCounter_231_reset = reset;
  assign SaturatingCounter_231_io_enable = _T_1037;
  assign SaturatingCounter_232_clock = clock;
  assign SaturatingCounter_232_reset = reset;
  assign SaturatingCounter_232_io_enable = _T_1038;
  assign SaturatingCounter_233_clock = clock;
  assign SaturatingCounter_233_reset = reset;
  assign SaturatingCounter_233_io_enable = _T_1044;
  assign SaturatingCounter_234_clock = clock;
  assign SaturatingCounter_234_reset = reset;
  assign SaturatingCounter_234_io_enable = _T_1045;
  assign SaturatingCounter_235_clock = clock;
  assign SaturatingCounter_235_reset = reset;
  assign SaturatingCounter_235_io_enable = _T_1051;
  assign SaturatingCounter_236_clock = clock;
  assign SaturatingCounter_236_reset = reset;
  assign SaturatingCounter_236_io_enable = _T_1052;
  assign SaturatingCounter_237_clock = clock;
  assign SaturatingCounter_237_reset = reset;
  assign SaturatingCounter_237_io_enable = _T_1058;
  assign SaturatingCounter_238_clock = clock;
  assign SaturatingCounter_238_reset = reset;
  assign SaturatingCounter_238_io_enable = _T_1059;
  assign SaturatingCounter_239_clock = clock;
  assign SaturatingCounter_239_reset = reset;
  assign SaturatingCounter_239_io_enable = _T_1065;
  assign SaturatingCounter_240_clock = clock;
  assign SaturatingCounter_240_reset = reset;
  assign SaturatingCounter_240_io_enable = _T_1066;
  assign SaturatingCounter_241_clock = clock;
  assign SaturatingCounter_241_reset = reset;
  assign SaturatingCounter_241_io_enable = _T_1072;
  assign SaturatingCounter_242_clock = clock;
  assign SaturatingCounter_242_reset = reset;
  assign SaturatingCounter_242_io_enable = _T_1073;
  assign SaturatingCounter_243_clock = clock;
  assign SaturatingCounter_243_reset = reset;
  assign SaturatingCounter_243_io_enable = _T_1079;
  assign SaturatingCounter_244_clock = clock;
  assign SaturatingCounter_244_reset = reset;
  assign SaturatingCounter_244_io_enable = _T_1080;
  assign SaturatingCounter_245_clock = clock;
  assign SaturatingCounter_245_reset = reset;
  assign SaturatingCounter_245_io_enable = _T_1086;
  assign SaturatingCounter_246_clock = clock;
  assign SaturatingCounter_246_reset = reset;
  assign SaturatingCounter_246_io_enable = _T_1087;
  assign SaturatingCounter_247_clock = clock;
  assign SaturatingCounter_247_reset = reset;
  assign SaturatingCounter_247_io_enable = _T_1093;
  assign SaturatingCounter_248_clock = clock;
  assign SaturatingCounter_248_reset = reset;
  assign SaturatingCounter_248_io_enable = _T_1094;
  assign SaturatingCounter_249_clock = clock;
  assign SaturatingCounter_249_reset = reset;
  assign SaturatingCounter_249_io_enable = _T_1100;
  assign SaturatingCounter_250_clock = clock;
  assign SaturatingCounter_250_reset = reset;
  assign SaturatingCounter_250_io_enable = _T_1101;
  assign SaturatingCounter_251_clock = clock;
  assign SaturatingCounter_251_reset = reset;
  assign SaturatingCounter_251_io_enable = _T_1107;
  assign SaturatingCounter_252_clock = clock;
  assign SaturatingCounter_252_reset = reset;
  assign SaturatingCounter_252_io_enable = _T_1108;
  assign SaturatingCounter_253_clock = clock;
  assign SaturatingCounter_253_reset = reset;
  assign SaturatingCounter_253_io_enable = _T_1114;
  assign SaturatingCounter_254_clock = clock;
  assign SaturatingCounter_254_reset = reset;
  assign SaturatingCounter_254_io_enable = _T_1115;
  assign SaturatingCounter_255_clock = clock;
  assign SaturatingCounter_255_reset = reset;
  assign SaturatingCounter_255_io_enable = _T_1121;
  assign SaturatingCounter_256_clock = clock;
  assign SaturatingCounter_256_reset = reset;
  assign SaturatingCounter_256_io_enable = _T_1122;
  assign SaturatingCounter_257_clock = clock;
  assign SaturatingCounter_257_reset = reset;
  assign SaturatingCounter_257_io_enable = _T_1128;
  assign SaturatingCounter_258_clock = clock;
  assign SaturatingCounter_258_reset = reset;
  assign SaturatingCounter_258_io_enable = _T_1129;
  assign SaturatingCounter_259_clock = clock;
  assign SaturatingCounter_259_reset = reset;
  assign SaturatingCounter_259_io_enable = _T_1135;
  assign SaturatingCounter_260_clock = clock;
  assign SaturatingCounter_260_reset = reset;
  assign SaturatingCounter_260_io_enable = _T_1136;
  assign SaturatingCounter_261_clock = clock;
  assign SaturatingCounter_261_reset = reset;
  assign SaturatingCounter_261_io_enable = _T_1142;
  assign SaturatingCounter_262_clock = clock;
  assign SaturatingCounter_262_reset = reset;
  assign SaturatingCounter_262_io_enable = _T_1143;
  assign SaturatingCounter_263_clock = clock;
  assign SaturatingCounter_263_reset = reset;
  assign SaturatingCounter_263_io_enable = _T_1149;
  assign SaturatingCounter_264_clock = clock;
  assign SaturatingCounter_264_reset = reset;
  assign SaturatingCounter_264_io_enable = _T_1150;
  assign SaturatingCounter_265_clock = clock;
  assign SaturatingCounter_265_reset = reset;
  assign SaturatingCounter_265_io_enable = _T_1156;
  assign SaturatingCounter_266_clock = clock;
  assign SaturatingCounter_266_reset = reset;
  assign SaturatingCounter_266_io_enable = _T_1157;
  assign SaturatingCounter_267_clock = clock;
  assign SaturatingCounter_267_reset = reset;
  assign SaturatingCounter_267_io_enable = _T_1163;
  assign SaturatingCounter_268_clock = clock;
  assign SaturatingCounter_268_reset = reset;
  assign SaturatingCounter_268_io_enable = _T_1164;
  assign SaturatingCounter_269_clock = clock;
  assign SaturatingCounter_269_reset = reset;
  assign SaturatingCounter_269_io_enable = _T_1170;
  assign SaturatingCounter_270_clock = clock;
  assign SaturatingCounter_270_reset = reset;
  assign SaturatingCounter_270_io_enable = _T_1171;
  assign SaturatingCounter_271_clock = clock;
  assign SaturatingCounter_271_reset = reset;
  assign SaturatingCounter_271_io_enable = _T_1177;
  assign SaturatingCounter_272_clock = clock;
  assign SaturatingCounter_272_reset = reset;
  assign SaturatingCounter_272_io_enable = _T_1178;
  assign SaturatingCounter_273_clock = clock;
  assign SaturatingCounter_273_reset = reset;
  assign SaturatingCounter_273_io_enable = _T_1184;
  assign SaturatingCounter_274_clock = clock;
  assign SaturatingCounter_274_reset = reset;
  assign SaturatingCounter_274_io_enable = _T_1185;
  assign SaturatingCounter_275_clock = clock;
  assign SaturatingCounter_275_reset = reset;
  assign SaturatingCounter_275_io_enable = _T_1191;
  assign SaturatingCounter_276_clock = clock;
  assign SaturatingCounter_276_reset = reset;
  assign SaturatingCounter_276_io_enable = _T_1192;
  assign SaturatingCounter_277_clock = clock;
  assign SaturatingCounter_277_reset = reset;
  assign SaturatingCounter_277_io_enable = _T_1198;
  assign SaturatingCounter_278_clock = clock;
  assign SaturatingCounter_278_reset = reset;
  assign SaturatingCounter_278_io_enable = _T_1199;
  assign SaturatingCounter_279_clock = clock;
  assign SaturatingCounter_279_reset = reset;
  assign SaturatingCounter_279_io_enable = _T_1205;
  assign SaturatingCounter_280_clock = clock;
  assign SaturatingCounter_280_reset = reset;
  assign SaturatingCounter_280_io_enable = _T_1206;
  assign SaturatingCounter_281_clock = clock;
  assign SaturatingCounter_281_reset = reset;
  assign SaturatingCounter_281_io_enable = _T_1212;
  assign SaturatingCounter_282_clock = clock;
  assign SaturatingCounter_282_reset = reset;
  assign SaturatingCounter_282_io_enable = _T_1213;
  assign SaturatingCounter_283_clock = clock;
  assign SaturatingCounter_283_reset = reset;
  assign SaturatingCounter_283_io_enable = _T_1219;
  assign SaturatingCounter_284_clock = clock;
  assign SaturatingCounter_284_reset = reset;
  assign SaturatingCounter_284_io_enable = _T_1220;
  assign SaturatingCounter_285_clock = clock;
  assign SaturatingCounter_285_reset = reset;
  assign SaturatingCounter_285_io_enable = _T_1226;
  assign SaturatingCounter_286_clock = clock;
  assign SaturatingCounter_286_reset = reset;
  assign SaturatingCounter_286_io_enable = _T_1227;
  assign SaturatingCounter_287_clock = clock;
  assign SaturatingCounter_287_reset = reset;
  assign SaturatingCounter_287_io_enable = _T_1233;
  assign SaturatingCounter_288_clock = clock;
  assign SaturatingCounter_288_reset = reset;
  assign SaturatingCounter_288_io_enable = _T_1234;
  assign SaturatingCounter_289_clock = clock;
  assign SaturatingCounter_289_reset = reset;
  assign SaturatingCounter_289_io_enable = _T_1240;
  assign SaturatingCounter_290_clock = clock;
  assign SaturatingCounter_290_reset = reset;
  assign SaturatingCounter_290_io_enable = _T_1241;
  assign SaturatingCounter_291_clock = clock;
  assign SaturatingCounter_291_reset = reset;
  assign SaturatingCounter_291_io_enable = _T_1247;
  assign SaturatingCounter_292_clock = clock;
  assign SaturatingCounter_292_reset = reset;
  assign SaturatingCounter_292_io_enable = _T_1248;
  assign SaturatingCounter_293_clock = clock;
  assign SaturatingCounter_293_reset = reset;
  assign SaturatingCounter_293_io_enable = _T_1254;
  assign SaturatingCounter_294_clock = clock;
  assign SaturatingCounter_294_reset = reset;
  assign SaturatingCounter_294_io_enable = _T_1255;
  assign SaturatingCounter_295_clock = clock;
  assign SaturatingCounter_295_reset = reset;
  assign SaturatingCounter_295_io_enable = _T_1261;
  assign SaturatingCounter_296_clock = clock;
  assign SaturatingCounter_296_reset = reset;
  assign SaturatingCounter_296_io_enable = _T_1262;
  assign SaturatingCounter_297_clock = clock;
  assign SaturatingCounter_297_reset = reset;
  assign SaturatingCounter_297_io_enable = _T_1268;
  assign SaturatingCounter_298_clock = clock;
  assign SaturatingCounter_298_reset = reset;
  assign SaturatingCounter_298_io_enable = _T_1269;
  assign SaturatingCounter_299_clock = clock;
  assign SaturatingCounter_299_reset = reset;
  assign SaturatingCounter_299_io_enable = _T_1275;
  assign SaturatingCounter_300_clock = clock;
  assign SaturatingCounter_300_reset = reset;
  assign SaturatingCounter_300_io_enable = _T_1276;
  assign SaturatingCounter_301_clock = clock;
  assign SaturatingCounter_301_reset = reset;
  assign SaturatingCounter_301_io_enable = _T_1282;
  assign SaturatingCounter_302_clock = clock;
  assign SaturatingCounter_302_reset = reset;
  assign SaturatingCounter_302_io_enable = _T_1283;
  assign SaturatingCounter_303_clock = clock;
  assign SaturatingCounter_303_reset = reset;
  assign SaturatingCounter_303_io_enable = _T_1289;
  assign SaturatingCounter_304_clock = clock;
  assign SaturatingCounter_304_reset = reset;
  assign SaturatingCounter_304_io_enable = _T_1290;
  assign SaturatingCounter_305_clock = clock;
  assign SaturatingCounter_305_reset = reset;
  assign SaturatingCounter_305_io_enable = _T_1296;
  assign SaturatingCounter_306_clock = clock;
  assign SaturatingCounter_306_reset = reset;
  assign SaturatingCounter_306_io_enable = _T_1297;
  assign SaturatingCounter_307_clock = clock;
  assign SaturatingCounter_307_reset = reset;
  assign SaturatingCounter_307_io_enable = _T_1303;
  assign SaturatingCounter_308_clock = clock;
  assign SaturatingCounter_308_reset = reset;
  assign SaturatingCounter_308_io_enable = _T_1304;
  assign SaturatingCounter_309_clock = clock;
  assign SaturatingCounter_309_reset = reset;
  assign SaturatingCounter_309_io_enable = _T_1310;
  assign SaturatingCounter_310_clock = clock;
  assign SaturatingCounter_310_reset = reset;
  assign SaturatingCounter_310_io_enable = _T_1311;
  assign SaturatingCounter_311_clock = clock;
  assign SaturatingCounter_311_reset = reset;
  assign SaturatingCounter_311_io_enable = _T_1317;
  assign SaturatingCounter_312_clock = clock;
  assign SaturatingCounter_312_reset = reset;
  assign SaturatingCounter_312_io_enable = _T_1318;
  assign SaturatingCounter_313_clock = clock;
  assign SaturatingCounter_313_reset = reset;
  assign SaturatingCounter_313_io_enable = _T_1324;
  assign SaturatingCounter_314_clock = clock;
  assign SaturatingCounter_314_reset = reset;
  assign SaturatingCounter_314_io_enable = _T_1325;
  assign SaturatingCounter_315_clock = clock;
  assign SaturatingCounter_315_reset = reset;
  assign SaturatingCounter_315_io_enable = _T_1331;
  assign SaturatingCounter_316_clock = clock;
  assign SaturatingCounter_316_reset = reset;
  assign SaturatingCounter_316_io_enable = _T_1332;
  assign SaturatingCounter_317_clock = clock;
  assign SaturatingCounter_317_reset = reset;
  assign SaturatingCounter_317_io_enable = _T_1338;
  assign SaturatingCounter_318_clock = clock;
  assign SaturatingCounter_318_reset = reset;
  assign SaturatingCounter_318_io_enable = _T_1339;
  assign SaturatingCounter_319_clock = clock;
  assign SaturatingCounter_319_reset = reset;
  assign SaturatingCounter_319_io_enable = _T_1345;
  assign SaturatingCounter_320_clock = clock;
  assign SaturatingCounter_320_reset = reset;
  assign SaturatingCounter_320_io_enable = _T_1346;
  assign SaturatingCounter_321_clock = clock;
  assign SaturatingCounter_321_reset = reset;
  assign SaturatingCounter_321_io_enable = _T_1352;
  assign SaturatingCounter_322_clock = clock;
  assign SaturatingCounter_322_reset = reset;
  assign SaturatingCounter_322_io_enable = _T_1353;
  assign SaturatingCounter_323_clock = clock;
  assign SaturatingCounter_323_reset = reset;
  assign SaturatingCounter_323_io_enable = _T_1359;
  assign SaturatingCounter_324_clock = clock;
  assign SaturatingCounter_324_reset = reset;
  assign SaturatingCounter_324_io_enable = _T_1360;
  assign SaturatingCounter_325_clock = clock;
  assign SaturatingCounter_325_reset = reset;
  assign SaturatingCounter_325_io_enable = _T_1366;
  assign SaturatingCounter_326_clock = clock;
  assign SaturatingCounter_326_reset = reset;
  assign SaturatingCounter_326_io_enable = _T_1367;
  assign SaturatingCounter_327_clock = clock;
  assign SaturatingCounter_327_reset = reset;
  assign SaturatingCounter_327_io_enable = _T_1373;
  assign SaturatingCounter_328_clock = clock;
  assign SaturatingCounter_328_reset = reset;
  assign SaturatingCounter_328_io_enable = _T_1374;
  assign SaturatingCounter_329_clock = clock;
  assign SaturatingCounter_329_reset = reset;
  assign SaturatingCounter_329_io_enable = _T_1380;
  assign SaturatingCounter_330_clock = clock;
  assign SaturatingCounter_330_reset = reset;
  assign SaturatingCounter_330_io_enable = _T_1381;
  assign SaturatingCounter_331_clock = clock;
  assign SaturatingCounter_331_reset = reset;
  assign SaturatingCounter_331_io_enable = _T_1387;
  assign SaturatingCounter_332_clock = clock;
  assign SaturatingCounter_332_reset = reset;
  assign SaturatingCounter_332_io_enable = _T_1388;
  assign SaturatingCounter_333_clock = clock;
  assign SaturatingCounter_333_reset = reset;
  assign SaturatingCounter_333_io_enable = _T_1394;
  assign SaturatingCounter_334_clock = clock;
  assign SaturatingCounter_334_reset = reset;
  assign SaturatingCounter_334_io_enable = _T_1395;
  assign SaturatingCounter_335_clock = clock;
  assign SaturatingCounter_335_reset = reset;
  assign SaturatingCounter_335_io_enable = _T_1401;
  assign SaturatingCounter_336_clock = clock;
  assign SaturatingCounter_336_reset = reset;
  assign SaturatingCounter_336_io_enable = _T_1402;
  assign SaturatingCounter_337_clock = clock;
  assign SaturatingCounter_337_reset = reset;
  assign SaturatingCounter_337_io_enable = _T_1408;
  assign SaturatingCounter_338_clock = clock;
  assign SaturatingCounter_338_reset = reset;
  assign SaturatingCounter_338_io_enable = _T_1409;
  assign SaturatingCounter_339_clock = clock;
  assign SaturatingCounter_339_reset = reset;
  assign SaturatingCounter_339_io_enable = _T_1415;
  assign SaturatingCounter_340_clock = clock;
  assign SaturatingCounter_340_reset = reset;
  assign SaturatingCounter_340_io_enable = _T_1416;
  assign SaturatingCounter_341_clock = clock;
  assign SaturatingCounter_341_reset = reset;
  assign SaturatingCounter_341_io_enable = _T_1422;
  assign SaturatingCounter_342_clock = clock;
  assign SaturatingCounter_342_reset = reset;
  assign SaturatingCounter_342_io_enable = _T_1423;
  assign SaturatingCounter_343_clock = clock;
  assign SaturatingCounter_343_reset = reset;
  assign SaturatingCounter_343_io_enable = _T_1429;
  assign SaturatingCounter_344_clock = clock;
  assign SaturatingCounter_344_reset = reset;
  assign SaturatingCounter_344_io_enable = _T_1430;
  assign SaturatingCounter_345_clock = clock;
  assign SaturatingCounter_345_reset = reset;
  assign SaturatingCounter_345_io_enable = _T_1436;
  assign SaturatingCounter_346_clock = clock;
  assign SaturatingCounter_346_reset = reset;
  assign SaturatingCounter_346_io_enable = _T_1437;
  assign SaturatingCounter_347_clock = clock;
  assign SaturatingCounter_347_reset = reset;
  assign SaturatingCounter_347_io_enable = _T_1443;
  assign SaturatingCounter_348_clock = clock;
  assign SaturatingCounter_348_reset = reset;
  assign SaturatingCounter_348_io_enable = _T_1444;
  assign SaturatingCounter_349_clock = clock;
  assign SaturatingCounter_349_reset = reset;
  assign SaturatingCounter_349_io_enable = _T_1450;
  assign SaturatingCounter_350_clock = clock;
  assign SaturatingCounter_350_reset = reset;
  assign SaturatingCounter_350_io_enable = _T_1451;
  assign SaturatingCounter_351_clock = clock;
  assign SaturatingCounter_351_reset = reset;
  assign SaturatingCounter_351_io_enable = _T_1457;
  assign SaturatingCounter_352_clock = clock;
  assign SaturatingCounter_352_reset = reset;
  assign SaturatingCounter_352_io_enable = _T_1458;
  assign SaturatingCounter_353_clock = clock;
  assign SaturatingCounter_353_reset = reset;
  assign SaturatingCounter_353_io_enable = _T_1464;
  assign SaturatingCounter_354_clock = clock;
  assign SaturatingCounter_354_reset = reset;
  assign SaturatingCounter_354_io_enable = _T_1465;
  assign SaturatingCounter_355_clock = clock;
  assign SaturatingCounter_355_reset = reset;
  assign SaturatingCounter_355_io_enable = _T_1471;
  assign SaturatingCounter_356_clock = clock;
  assign SaturatingCounter_356_reset = reset;
  assign SaturatingCounter_356_io_enable = _T_1472;
  assign SaturatingCounter_357_clock = clock;
  assign SaturatingCounter_357_reset = reset;
  assign SaturatingCounter_357_io_enable = _T_1478;
  assign SaturatingCounter_358_clock = clock;
  assign SaturatingCounter_358_reset = reset;
  assign SaturatingCounter_358_io_enable = _T_1479;
  assign SaturatingCounter_359_clock = clock;
  assign SaturatingCounter_359_reset = reset;
  assign SaturatingCounter_359_io_enable = _T_1485;
  assign SaturatingCounter_360_clock = clock;
  assign SaturatingCounter_360_reset = reset;
  assign SaturatingCounter_360_io_enable = _T_1486;
  assign SaturatingCounter_361_clock = clock;
  assign SaturatingCounter_361_reset = reset;
  assign SaturatingCounter_361_io_enable = _T_1492;
  assign SaturatingCounter_362_clock = clock;
  assign SaturatingCounter_362_reset = reset;
  assign SaturatingCounter_362_io_enable = _T_1493;
  assign SaturatingCounter_363_clock = clock;
  assign SaturatingCounter_363_reset = reset;
  assign SaturatingCounter_363_io_enable = _T_1499;
  assign SaturatingCounter_364_clock = clock;
  assign SaturatingCounter_364_reset = reset;
  assign SaturatingCounter_364_io_enable = _T_1500;
  assign SaturatingCounter_365_clock = clock;
  assign SaturatingCounter_365_reset = reset;
  assign SaturatingCounter_365_io_enable = _T_1506;
  assign SaturatingCounter_366_clock = clock;
  assign SaturatingCounter_366_reset = reset;
  assign SaturatingCounter_366_io_enable = _T_1507;
  assign SaturatingCounter_367_clock = clock;
  assign SaturatingCounter_367_reset = reset;
  assign SaturatingCounter_367_io_enable = _T_1513;
  assign SaturatingCounter_368_clock = clock;
  assign SaturatingCounter_368_reset = reset;
  assign SaturatingCounter_368_io_enable = _T_1514;
  assign SaturatingCounter_369_clock = clock;
  assign SaturatingCounter_369_reset = reset;
  assign SaturatingCounter_369_io_enable = _T_1520;
  assign SaturatingCounter_370_clock = clock;
  assign SaturatingCounter_370_reset = reset;
  assign SaturatingCounter_370_io_enable = _T_1521;
  assign SaturatingCounter_371_clock = clock;
  assign SaturatingCounter_371_reset = reset;
  assign SaturatingCounter_371_io_enable = _T_1527;
  assign SaturatingCounter_372_clock = clock;
  assign SaturatingCounter_372_reset = reset;
  assign SaturatingCounter_372_io_enable = _T_1528;
  assign SaturatingCounter_373_clock = clock;
  assign SaturatingCounter_373_reset = reset;
  assign SaturatingCounter_373_io_enable = _T_1534;
  assign SaturatingCounter_374_clock = clock;
  assign SaturatingCounter_374_reset = reset;
  assign SaturatingCounter_374_io_enable = _T_1535;
  assign SaturatingCounter_375_clock = clock;
  assign SaturatingCounter_375_reset = reset;
  assign SaturatingCounter_375_io_enable = _T_1541;
  assign SaturatingCounter_376_clock = clock;
  assign SaturatingCounter_376_reset = reset;
  assign SaturatingCounter_376_io_enable = _T_1542;
  assign SaturatingCounter_377_clock = clock;
  assign SaturatingCounter_377_reset = reset;
  assign SaturatingCounter_377_io_enable = _T_1548;
  assign SaturatingCounter_378_clock = clock;
  assign SaturatingCounter_378_reset = reset;
  assign SaturatingCounter_378_io_enable = _T_1549;
  assign SaturatingCounter_379_clock = clock;
  assign SaturatingCounter_379_reset = reset;
  assign SaturatingCounter_379_io_enable = _T_1555;
  assign SaturatingCounter_380_clock = clock;
  assign SaturatingCounter_380_reset = reset;
  assign SaturatingCounter_380_io_enable = _T_1556;
  assign SaturatingCounter_381_clock = clock;
  assign SaturatingCounter_381_reset = reset;
  assign SaturatingCounter_381_io_enable = _T_1562;
  assign SaturatingCounter_382_clock = clock;
  assign SaturatingCounter_382_reset = reset;
  assign SaturatingCounter_382_io_enable = _T_1563;
endmodule
