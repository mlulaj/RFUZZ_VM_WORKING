module Sodor3Stage( // @[:Sodor3Stage.fir@3963.2]
  input          metaReset,
  input          clock, // @[:Sodor3Stage.fir@3964.4]
  input          reset, // @[:Sodor3Stage.fir@3965.4]
  input          io_imem_req_ready, // @[:Sodor3Stage.fir@3966.4]
  output         io_imem_req_valid, // @[:Sodor3Stage.fir@3966.4]
  output [31:0]  io_imem_req_bits_addr, // @[:Sodor3Stage.fir@3966.4]
  output [31:0]  io_imem_req_bits_data, // @[:Sodor3Stage.fir@3966.4]
  output         io_imem_req_bits_fcn, // @[:Sodor3Stage.fir@3966.4]
  output [2:0]   io_imem_req_bits_typ, // @[:Sodor3Stage.fir@3966.4]
  input          io_imem_resp_valid, // @[:Sodor3Stage.fir@3966.4]
  input  [31:0]  io_imem_resp_bits_data, // @[:Sodor3Stage.fir@3966.4]
  input          io_reset, // @[:Sodor3Stage.fir@3966.4]
  output         assert_out,
  output [745:0] auto_cover_out
);
  wire  core_metaReset; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core_clock; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core_reset; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire [31:0] core_io_imem_req_bits_addr; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire [31:0] core_io_imem_resp_bits_data; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire [31:0] core_io_dmem_req_bits_addr; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire [31:0] core_io_dmem_req_bits_data; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core_io_dmem_req_bits_fcn; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire [2:0] core_io_dmem_req_bits_typ; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire [31:0] core_io_dmem_resp_bits_data; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_338; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_224; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_218; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_21; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_91; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_323; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_302; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_51; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_304; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_199; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_6; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_148; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_239; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_403; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_1; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_24; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_247; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_106; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_317; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_133; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_205; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_385; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_39; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_232; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_418; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_127; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_197; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_331; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_190; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_12; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_226; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_296; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_9_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_45; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_112; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_298; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_203; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_72; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_211; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_325; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_397; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_424; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_30; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_310; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_319; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_66; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_9_1; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_212; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_220; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_214; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_100; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_109; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_320; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_313; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_282; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_200; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_177; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_208; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_388; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_391; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_381; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_412; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_27; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_276; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_191; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_181; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_54; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_193; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_190_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_15; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_289; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_12_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_406; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_299; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_48; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_115; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_311; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_206; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_367; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_175; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_6_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_305; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_33; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_274; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_121; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_307; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_373; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_375; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_229; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_94; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_292; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_183; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_376; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_382; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_0_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_10; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_370; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_349; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_196; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_186; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_262; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_400; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_103; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_264; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_295; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_355; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_159; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_202; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_171; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_357; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_270; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_277; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_384; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_36; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_285; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_165; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_279; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_194; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_184; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_378; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_293; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_21_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_301; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_157; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_3_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_361; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_394; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_15_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_256; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_363; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_9_2; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_258; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_97; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_283; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_163; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_178; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_345; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_339; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_8; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_11; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_18; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_259; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_147; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_358; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_330; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_172; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_86; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_13; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_271; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_265; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_280; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_160; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_273; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_343; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_379; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_351; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_238; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_231; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_189; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_337; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_153; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_288; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_364; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_244; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_366; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_252; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_180; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_166; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_71; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_174; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_168; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_372; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_3_1; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_387; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_246; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_267; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_286; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_151; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_187; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_354; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_213; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_249; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_319_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_268; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_240; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_141; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_135; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_226_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_234; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_348; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_261; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_312; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_53; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_333; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_147_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_68; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_156; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_352; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_247_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_360; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_369; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_325_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_2; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_74; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_327; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_169; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_89; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_162; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_232_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_426; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_7_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_331_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_129; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_346; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_154; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_340; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_253; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_228; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_411; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_255; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_120; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_211_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_80; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_220_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_342; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_229_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_393; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_292_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_307_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_193_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_56; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_144; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_17; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_11_1; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_408; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_222; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_313_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_117; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_328; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_321; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_2_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_235; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_243; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_237; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_123; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_102; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_3_2; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_62; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_150; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_336; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_201; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_195; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_23; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_414; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_250; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_300; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_294; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_309; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_77; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_208_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_83; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_214_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_216; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_241; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_420; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_35; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_5_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_41; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_315; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_429; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_138; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_334; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_217; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_402; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_17_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_225; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_105; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_316; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_50; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_44; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_324; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_180_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_318; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_384_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_396; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_386; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_38; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_301_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_196_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_186_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_65; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_295_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_20; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_223; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_23_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_417; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_111; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_322; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_210; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_5_1; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_219; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_279_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_310_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_285_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_423; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_132; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_126; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_287; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_202_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_378_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_90; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_204; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_99; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_303; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_297; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_59; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_188; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_198; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_351_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_176; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_387_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_11_2; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_380; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_93; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_161; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_192; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_189_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_14_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_372_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_207; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_267_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_405; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_260; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_26; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_114; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_269; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_174_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_205_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_182; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_399; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_368; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_273_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_390; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_32; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_281; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_275; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_291; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_168_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_47; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_199_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_5_2; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_389; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_298_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_304_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_306; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_366_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_8_1; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_374; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_108; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_360_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_288_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_356; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_375_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_255_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_261_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_20_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_14_1; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_29; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_270_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_150_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_333_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_82; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_177_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_170; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_381_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_185; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_1_1; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_276_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_10_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_278; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_143; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_354_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_348_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_249_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_96; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_9_3; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_263; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_164; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_158; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_369_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_183_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_362; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_377; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_257; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_282_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_284; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_179; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_383; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_242; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_8_2; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_162_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_156_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_341; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_76; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_165_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_173; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_224_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_359; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_251; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_131; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_7_1; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_146; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_342_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_350; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_344; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_239_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_264_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_272; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_64; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_58; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_159_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_222_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_363_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_357_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_230; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_365; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_321_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_7_2; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_330_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_323_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_85; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_338_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_79; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_243_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_2_2; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_237_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_245; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_12_1; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_315_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_336_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_70; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_152; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_167; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_422; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_258_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_371; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_266; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_125; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_171_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_212_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_303_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_254; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_146_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_13_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_155; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_149; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_225_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_227; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_113; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_140; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_326; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_7_3; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_231_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_425; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_404; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_240_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_353; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_248; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_107; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_6_3; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_311_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_339_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_153_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_73; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_67; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_347; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_206_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_252_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_410; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_297_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_419; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_233; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_305_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_128; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_324_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_332; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_219_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_88; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_1_3; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_246_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_318_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_52; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_46; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_134; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_345_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_204_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_213_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_228_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_221; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_407; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_382_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_28; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_281_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_4_1; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_40; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_55; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_329; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_194_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_392; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_0_2; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_234_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_10_2; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_236; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_101; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_312_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_192_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_306_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_61; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_207_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_16; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_22; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_300_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_34; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_116; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_122; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_327_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_182_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_320_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_215; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_335; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_291_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_290; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_293_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_428; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_49; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_137; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_200_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_209; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_95; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_413; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_314; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_308; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_4_2; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_383_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_16_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_395; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_385_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_104; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_195_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_302_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_317_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_203_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_172_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_197_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_370_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_416; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_22_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_271_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_119; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_185_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_179_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_216_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_379_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_187_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_401; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_43; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_278_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_296_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_286_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_201_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_364_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_1_4; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_210_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_98; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_263_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_309_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_37; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_164_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_110; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_362_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_19; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_377_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_218_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_294_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_284_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_371_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_260_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_266_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_380_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_25; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_365_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_181_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_175_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_251_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_15_1; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_289_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_359_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_352_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_14_2; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_152_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_31; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_274_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_160_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_169_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_191_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_188_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_373_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_19_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_367_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_268_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_173_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_290_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_280_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_287_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_154_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_87; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_299_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_386_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_10_3; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_245_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_398; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_4_3; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_388_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_253_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_92; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_5_3; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_272_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_344_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_198_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_167_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_346_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_334_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_340_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_254_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_13_2; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_3_4; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_256_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_328_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_161_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_347_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_81; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_355_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_170_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_7_5; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_8_3; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_275_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_269_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_155_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_277_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_69; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_157_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_368_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_233_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_227_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_235_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_184_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_326_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_149_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_60; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_283_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_142; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_353_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_178_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_248_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_241_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_361_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_136; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_75; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_163_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_349_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_374_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_427; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_376_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_262_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_332_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_176_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_166_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_358_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_314_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_308_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_42; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_265_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_316_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_130; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_124; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_341_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_343_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_223_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_238_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_118; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_5_4; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_151_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_145; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_337_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_18_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_356_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_244_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_409; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_11_3; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_322_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_158_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_209_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_78; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_217_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_221_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_236_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_421; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_415; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_335_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_329_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_63; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_230_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_242_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_257_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_6_4; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_57; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_250_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_259_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_139; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_350_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_215_0; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  core__GEN_84; // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
  wire  memory_metaReset; // @[top.scala 29:28:Sodor3Stage.fir@3974.4]
  wire  memory_clock; // @[top.scala 29:28:Sodor3Stage.fir@3974.4]
  wire [31:0] memory_io_core_ports_0_req_bits_addr; // @[top.scala 29:28:Sodor3Stage.fir@3974.4]
  wire [31:0] memory_io_core_ports_0_req_bits_data; // @[top.scala 29:28:Sodor3Stage.fir@3974.4]
  wire  memory_io_core_ports_0_req_bits_fcn; // @[top.scala 29:28:Sodor3Stage.fir@3974.4]
  wire [2:0] memory_io_core_ports_0_req_bits_typ; // @[top.scala 29:28:Sodor3Stage.fir@3974.4]
  wire [31:0] memory_io_core_ports_0_resp_bits_data; // @[top.scala 29:28:Sodor3Stage.fir@3974.4]
  wire  memory__GEN_3_0; // @[top.scala 29:28:Sodor3Stage.fir@3974.4]
  wire  memory__GEN_7_0; // @[top.scala 29:28:Sodor3Stage.fir@3974.4]
  wire  memory__GEN_1_1; // @[top.scala 29:28:Sodor3Stage.fir@3974.4]
  wire  memory__GEN_4_0; // @[top.scala 29:28:Sodor3Stage.fir@3974.4]
  wire  memory__GEN_2_2; // @[top.scala 29:28:Sodor3Stage.fir@3974.4]
  wire  memory__GEN_3_4; // @[top.scala 29:28:Sodor3Stage.fir@3974.4]
  wire  memory__GEN_6_3; // @[top.scala 29:28:Sodor3Stage.fir@3974.4]
  wire  memory__GEN_0_2; // @[top.scala 29:28:Sodor3Stage.fir@3974.4]
  wire  memory__GEN_1_3; // @[top.scala 29:28:Sodor3Stage.fir@3974.4]
  wire  memory__GEN_2_4; // @[top.scala 29:28:Sodor3Stage.fir@3974.4]
  wire  memory__GEN_0_4; // @[top.scala 29:28:Sodor3Stage.fir@3974.4]
  wire  memory__GEN_5_6; // @[top.scala 29:28:Sodor3Stage.fir@3974.4]
  wire  profilePin;
  wire  profilePin_0;
  wire [1:0] _GEN_749; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_1;
  wire [2:0] _GEN_750; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_2;
  wire [3:0] _GEN_751; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_3;
  wire [4:0] _GEN_752; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_4;
  wire [5:0] _GEN_753; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_5;
  wire [6:0] _GEN_754; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_6;
  wire [7:0] _GEN_755; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_7;
  wire [8:0] _GEN_756; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_8;
  wire [9:0] _GEN_757; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_9;
  wire [10:0] _GEN_758; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_10;
  wire [11:0] _GEN_759; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_11;
  wire [12:0] _GEN_760; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_12;
  wire [13:0] _GEN_761; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_13;
  wire [14:0] _GEN_762; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_14;
  wire [15:0] _GEN_763; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_15;
  wire [16:0] _GEN_764; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_16;
  wire [17:0] _GEN_765; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_17;
  wire [18:0] _GEN_766; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_18;
  wire [19:0] _GEN_767; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_19;
  wire [20:0] _GEN_768; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_20;
  wire [21:0] _GEN_769; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_21;
  wire [22:0] _GEN_770; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_22;
  wire [23:0] _GEN_771; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_23;
  wire [24:0] _GEN_772; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_24;
  wire [25:0] _GEN_773; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_25;
  wire [26:0] _GEN_774; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_26;
  wire [27:0] _GEN_775; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_27;
  wire [28:0] _GEN_776; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_28;
  wire [29:0] _GEN_777; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_29;
  wire [30:0] _GEN_778; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_30;
  wire [31:0] _GEN_779; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_31;
  wire [32:0] _GEN_780; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_32;
  wire [33:0] _GEN_781; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_33;
  wire [34:0] _GEN_782; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_34;
  wire [35:0] _GEN_783; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_35;
  wire [36:0] _GEN_784; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_36;
  wire [37:0] _GEN_785; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_37;
  wire [38:0] _GEN_786; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_38;
  wire [39:0] _GEN_787; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_39;
  wire [40:0] _GEN_788; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_40;
  wire [41:0] _GEN_789; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_41;
  wire [42:0] _GEN_790; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_42;
  wire [43:0] _GEN_791; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_43;
  wire [44:0] _GEN_792; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_44;
  wire [45:0] _GEN_793; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_45;
  wire [46:0] _GEN_794; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_46;
  wire [47:0] _GEN_795; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_47;
  wire [48:0] _GEN_796; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_48;
  wire [49:0] _GEN_797; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_49;
  wire [50:0] _GEN_798; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_50;
  wire [51:0] _GEN_799; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_51;
  wire [52:0] _GEN_800; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_52;
  wire [53:0] _GEN_801; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_53;
  wire [54:0] _GEN_802; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_54;
  wire [55:0] _GEN_803; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_55;
  wire [56:0] _GEN_804; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_56;
  wire [57:0] _GEN_805; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_57;
  wire [58:0] _GEN_806; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_58;
  wire [59:0] _GEN_807; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_59;
  wire [60:0] _GEN_808; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_60;
  wire [61:0] _GEN_809; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_61;
  wire [62:0] _GEN_810; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_62;
  wire [63:0] _GEN_811; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_63;
  wire [64:0] _GEN_812; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_64;
  wire [65:0] _GEN_813; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_65;
  wire [66:0] _GEN_814; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_66;
  wire [67:0] _GEN_815; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_67;
  wire [68:0] _GEN_816; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_68;
  wire [69:0] _GEN_817; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_69;
  wire [70:0] _GEN_818; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_70;
  wire [71:0] _GEN_819; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_71;
  wire [72:0] _GEN_820; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_72;
  wire [73:0] _GEN_821; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_73;
  wire [74:0] _GEN_822; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_74;
  wire [75:0] _GEN_823; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_75;
  wire [76:0] _GEN_824; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_76;
  wire [77:0] _GEN_825; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_77;
  wire [78:0] _GEN_826; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_78;
  wire [79:0] _GEN_827; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_79;
  wire [80:0] _GEN_828; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_80;
  wire [81:0] _GEN_829; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_81;
  wire [82:0] _GEN_830; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_82;
  wire [83:0] _GEN_831; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_83;
  wire [84:0] _GEN_832; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_84;
  wire [85:0] _GEN_833; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_85;
  wire [86:0] _GEN_834; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_86;
  wire [87:0] _GEN_835; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_87;
  wire [88:0] _GEN_836; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_88;
  wire [89:0] _GEN_837; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_89;
  wire [90:0] _GEN_838; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_90;
  wire [91:0] _GEN_839; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_91;
  wire [92:0] _GEN_840; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_92;
  wire [93:0] _GEN_841; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_93;
  wire [94:0] _GEN_842; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_94;
  wire [95:0] _GEN_843; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_95;
  wire [96:0] _GEN_844; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_96;
  wire [97:0] _GEN_845; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_97;
  wire [98:0] _GEN_846; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_98;
  wire [99:0] _GEN_847; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_99;
  wire [100:0] _GEN_848; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_100;
  wire [101:0] _GEN_849; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_101;
  wire [102:0] _GEN_850; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_102;
  wire [103:0] _GEN_851; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_103;
  wire [104:0] _GEN_852; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_104;
  wire [105:0] _GEN_853; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_105;
  wire [106:0] _GEN_854; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_106;
  wire [107:0] _GEN_855; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_107;
  wire [108:0] _GEN_856; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_108;
  wire [109:0] _GEN_857; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_109;
  wire [110:0] _GEN_858; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_110;
  wire [111:0] _GEN_859; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_111;
  wire [112:0] _GEN_860; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_112;
  wire [113:0] _GEN_861; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_113;
  wire [114:0] _GEN_862; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_114;
  wire [115:0] _GEN_863; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_115;
  wire [116:0] _GEN_864; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_116;
  wire [117:0] _GEN_865; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_117;
  wire [118:0] _GEN_866; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_118;
  wire [119:0] _GEN_867; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_119;
  wire [120:0] _GEN_868; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_120;
  wire [121:0] _GEN_869; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_121;
  wire [122:0] _GEN_870; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_122;
  wire [123:0] _GEN_871; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_123;
  wire [124:0] _GEN_872; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_124;
  wire [125:0] _GEN_873; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_125;
  wire [126:0] _GEN_874; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_126;
  wire [127:0] _GEN_875; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_127;
  wire [128:0] _GEN_876; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_128;
  wire [129:0] _GEN_877; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_129;
  wire [130:0] _GEN_878; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_130;
  wire [131:0] _GEN_879; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_131;
  wire [132:0] _GEN_880; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_132;
  wire [133:0] _GEN_881; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_133;
  wire [134:0] _GEN_882; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_134;
  wire [135:0] _GEN_883; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_135;
  wire [136:0] _GEN_884; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_136;
  wire [137:0] _GEN_885; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_137;
  wire [138:0] _GEN_886; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_138;
  wire [139:0] _GEN_887; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_139;
  wire [140:0] _GEN_888; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_140;
  wire [141:0] _GEN_889; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_141;
  wire [142:0] _GEN_890; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_142;
  wire [143:0] _GEN_891; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_143;
  wire [144:0] _GEN_892; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_144;
  wire [145:0] _GEN_893; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_145;
  wire [146:0] _GEN_894; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_146;
  wire [147:0] _GEN_895; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_147;
  wire [148:0] _GEN_896; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_148;
  wire [149:0] _GEN_897; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_149;
  wire [150:0] _GEN_898; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_150;
  wire [151:0] _GEN_899; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_151;
  wire [152:0] _GEN_900; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_152;
  wire [153:0] _GEN_901; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_153;
  wire [154:0] _GEN_902; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_154;
  wire [155:0] _GEN_903; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_155;
  wire [156:0] _GEN_904; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_156;
  wire [157:0] _GEN_905; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_157;
  wire [158:0] _GEN_906; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_158;
  wire [159:0] _GEN_907; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_159;
  wire [160:0] _GEN_908; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_160;
  wire [161:0] _GEN_909; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_161;
  wire [162:0] _GEN_910; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_162;
  wire [163:0] _GEN_911; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_163;
  wire [164:0] _GEN_912; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_164;
  wire [165:0] _GEN_913; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_165;
  wire [166:0] _GEN_914; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_166;
  wire [167:0] _GEN_915; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_167;
  wire [168:0] _GEN_916; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_168;
  wire [169:0] _GEN_917; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_169;
  wire [170:0] _GEN_918; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_170;
  wire [171:0] _GEN_919; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_171;
  wire [172:0] _GEN_920; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_172;
  wire [173:0] _GEN_921; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_173;
  wire [174:0] _GEN_922; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_174;
  wire [175:0] _GEN_923; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_175;
  wire [176:0] _GEN_924; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_176;
  wire [177:0] _GEN_925; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_177;
  wire [178:0] _GEN_926; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_178;
  wire [179:0] _GEN_927; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_179;
  wire [180:0] _GEN_928; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_180;
  wire [181:0] _GEN_929; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_181;
  wire [182:0] _GEN_930; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_182;
  wire [183:0] _GEN_931; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_183;
  wire [184:0] _GEN_932; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_184;
  wire [185:0] _GEN_933; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_185;
  wire [186:0] _GEN_934; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_186;
  wire [187:0] _GEN_935; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_187;
  wire [188:0] _GEN_936; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_188;
  wire [189:0] _GEN_937; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_189;
  wire [190:0] _GEN_938; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_190;
  wire [191:0] _GEN_939; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_191;
  wire [192:0] _GEN_940; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_192;
  wire [193:0] _GEN_941; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_193;
  wire [194:0] _GEN_942; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_194;
  wire [195:0] _GEN_943; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_195;
  wire [196:0] _GEN_944; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_196;
  wire [197:0] _GEN_945; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_197;
  wire [198:0] _GEN_946; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_198;
  wire [199:0] _GEN_947; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_199;
  wire [200:0] _GEN_948; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_200;
  wire [201:0] _GEN_949; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_201;
  wire [202:0] _GEN_950; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_202;
  wire [203:0] _GEN_951; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_203;
  wire [204:0] _GEN_952; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_204;
  wire [205:0] _GEN_953; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_205;
  wire [206:0] _GEN_954; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_206;
  wire [207:0] _GEN_955; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_207;
  wire [208:0] _GEN_956; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_208;
  wire [209:0] _GEN_957; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_209;
  wire [210:0] _GEN_958; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_210;
  wire [211:0] _GEN_959; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_211;
  wire [212:0] _GEN_960; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_212;
  wire [213:0] _GEN_961; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_213;
  wire [214:0] _GEN_962; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_214;
  wire [215:0] _GEN_963; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_215;
  wire [216:0] _GEN_964; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_216;
  wire [217:0] _GEN_965; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_217;
  wire [218:0] _GEN_966; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_218;
  wire [219:0] _GEN_967; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_219;
  wire [220:0] _GEN_968; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_220;
  wire [221:0] _GEN_969; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_221;
  wire [222:0] _GEN_970; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_222;
  wire [223:0] _GEN_971; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_223;
  wire [224:0] _GEN_972; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_224;
  wire [225:0] _GEN_973; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_225;
  wire [226:0] _GEN_974; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_226;
  wire [227:0] _GEN_975; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_227;
  wire [228:0] _GEN_976; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_228;
  wire [229:0] _GEN_977; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_229;
  wire [230:0] _GEN_978; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_230;
  wire [231:0] _GEN_979; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_231;
  wire [232:0] _GEN_980; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_232;
  wire [233:0] _GEN_981; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_233;
  wire [234:0] _GEN_982; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_234;
  wire [235:0] _GEN_983; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_235;
  wire [236:0] _GEN_984; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_236;
  wire [237:0] _GEN_985; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_237;
  wire [238:0] _GEN_986; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_238;
  wire [239:0] _GEN_987; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_239;
  wire [240:0] _GEN_988; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_240;
  wire [241:0] _GEN_989; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_241;
  wire [242:0] _GEN_990; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_242;
  wire [243:0] _GEN_991; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_243;
  wire [244:0] _GEN_992; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_244;
  wire [245:0] _GEN_993; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_245;
  wire [246:0] _GEN_994; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_246;
  wire [247:0] _GEN_995; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_247;
  wire [248:0] _GEN_996; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_248;
  wire [249:0] _GEN_997; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_249;
  wire [250:0] _GEN_998; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_250;
  wire [251:0] _GEN_999; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_251;
  wire [252:0] _GEN_1000; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_252;
  wire [253:0] _GEN_1001; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_253;
  wire [254:0] _GEN_1002; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_254;
  wire [255:0] _GEN_1003; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_255;
  wire [256:0] _GEN_1004; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_256;
  wire [257:0] _GEN_1005; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_257;
  wire [258:0] _GEN_1006; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_258;
  wire [259:0] _GEN_1007; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_259;
  wire [260:0] _GEN_1008; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_260;
  wire [261:0] _GEN_1009; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_261;
  wire [262:0] _GEN_1010; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_262;
  wire [263:0] _GEN_1011; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_263;
  wire [264:0] _GEN_1012; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_264;
  wire [265:0] _GEN_1013; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_265;
  wire [266:0] _GEN_1014; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_266;
  wire [267:0] _GEN_1015; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_267;
  wire [268:0] _GEN_1016; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_268;
  wire [269:0] _GEN_1017; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_269;
  wire [270:0] _GEN_1018; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_270;
  wire [271:0] _GEN_1019; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_271;
  wire [272:0] _GEN_1020; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_272;
  wire [273:0] _GEN_1021; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_273;
  wire [274:0] _GEN_1022; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_274;
  wire [275:0] _GEN_1023; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_275;
  wire [276:0] _GEN_1024; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_276;
  wire [277:0] _GEN_1025; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_277;
  wire [278:0] _GEN_1026; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_278;
  wire [279:0] _GEN_1027; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_279;
  wire [280:0] _GEN_1028; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_280;
  wire [281:0] _GEN_1029; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_281;
  wire [282:0] _GEN_1030; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_282;
  wire [283:0] _GEN_1031; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_283;
  wire [284:0] _GEN_1032; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_284;
  wire [285:0] _GEN_1033; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_285;
  wire [286:0] _GEN_1034; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_286;
  wire [287:0] _GEN_1035; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_287;
  wire [288:0] _GEN_1036; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_288;
  wire [289:0] _GEN_1037; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_289;
  wire [290:0] _GEN_1038; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_290;
  wire [291:0] _GEN_1039; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_291;
  wire [292:0] _GEN_1040; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_292;
  wire [293:0] _GEN_1041; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_293;
  wire [294:0] _GEN_1042; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_294;
  wire [295:0] _GEN_1043; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_295;
  wire [296:0] _GEN_1044; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_296;
  wire [297:0] _GEN_1045; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_297;
  wire [298:0] _GEN_1046; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_298;
  wire [299:0] _GEN_1047; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_299;
  wire [300:0] _GEN_1048; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_300;
  wire [301:0] _GEN_1049; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_301;
  wire [302:0] _GEN_1050; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_302;
  wire [303:0] _GEN_1051; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_303;
  wire [304:0] _GEN_1052; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_304;
  wire [305:0] _GEN_1053; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_305;
  wire [306:0] _GEN_1054; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_306;
  wire [307:0] _GEN_1055; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_307;
  wire [308:0] _GEN_1056; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_308;
  wire [309:0] _GEN_1057; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_309;
  wire [310:0] _GEN_1058; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_310;
  wire [311:0] _GEN_1059; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_311;
  wire [312:0] _GEN_1060; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_312;
  wire [313:0] _GEN_1061; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_313;
  wire [314:0] _GEN_1062; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_314;
  wire [315:0] _GEN_1063; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_315;
  wire [316:0] _GEN_1064; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_316;
  wire [317:0] _GEN_1065; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_317;
  wire [318:0] _GEN_1066; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_318;
  wire [319:0] _GEN_1067; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_319;
  wire [320:0] _GEN_1068; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_320;
  wire [321:0] _GEN_1069; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_321;
  wire [322:0] _GEN_1070; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_322;
  wire [323:0] _GEN_1071; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_323;
  wire [324:0] _GEN_1072; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_324;
  wire [325:0] _GEN_1073; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_325;
  wire [326:0] _GEN_1074; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_326;
  wire [327:0] _GEN_1075; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_327;
  wire [328:0] _GEN_1076; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_328;
  wire [329:0] _GEN_1077; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_329;
  wire [330:0] _GEN_1078; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_330;
  wire [331:0] _GEN_1079; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_331;
  wire [332:0] _GEN_1080; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_332;
  wire [333:0] _GEN_1081; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_333;
  wire [334:0] _GEN_1082; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_334;
  wire [335:0] _GEN_1083; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_335;
  wire [336:0] _GEN_1084; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_336;
  wire [337:0] _GEN_1085; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_337;
  wire [338:0] _GEN_1086; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_338;
  wire [339:0] _GEN_1087; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_339;
  wire [340:0] _GEN_1088; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_340;
  wire [341:0] _GEN_1089; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_341;
  wire [342:0] _GEN_1090; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_342;
  wire [343:0] _GEN_1091; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_343;
  wire [344:0] _GEN_1092; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_344;
  wire [345:0] _GEN_1093; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_345;
  wire [346:0] _GEN_1094; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_346;
  wire [347:0] _GEN_1095; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_347;
  wire [348:0] _GEN_1096; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_348;
  wire [349:0] _GEN_1097; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_349;
  wire [350:0] _GEN_1098; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_350;
  wire [351:0] _GEN_1099; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_351;
  wire [352:0] _GEN_1100; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_352;
  wire [353:0] _GEN_1101; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_353;
  wire [354:0] _GEN_1102; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_354;
  wire [355:0] _GEN_1103; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_355;
  wire [356:0] _GEN_1104; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_356;
  wire [357:0] _GEN_1105; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_357;
  wire [358:0] _GEN_1106; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_358;
  wire [359:0] _GEN_1107; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_359;
  wire [360:0] _GEN_1108; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_360;
  wire [361:0] _GEN_1109; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_361;
  wire [362:0] _GEN_1110; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_362;
  wire [363:0] _GEN_1111; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_363;
  wire [364:0] _GEN_1112; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_364;
  wire [365:0] _GEN_1113; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_365;
  wire [366:0] _GEN_1114; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_366;
  wire [367:0] _GEN_1115; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_367;
  wire [368:0] _GEN_1116; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_368;
  wire [369:0] _GEN_1117; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_369;
  wire [370:0] _GEN_1118; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_370;
  wire [371:0] _GEN_1119; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_371;
  wire [372:0] _GEN_1120; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_372;
  wire [373:0] _GEN_1121; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_373;
  wire [374:0] _GEN_1122; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_374;
  wire [375:0] _GEN_1123; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_375;
  wire [376:0] _GEN_1124; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_376;
  wire [377:0] _GEN_1125; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_377;
  wire [378:0] _GEN_1126; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_378;
  wire [379:0] _GEN_1127; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_379;
  wire [380:0] _GEN_1128; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_380;
  wire [381:0] _GEN_1129; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_381;
  wire [382:0] _GEN_1130; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_382;
  wire [383:0] _GEN_1131; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_383;
  wire [384:0] _GEN_1132; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_384;
  wire [385:0] _GEN_1133; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_385;
  wire [386:0] _GEN_1134; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_386;
  wire [387:0] _GEN_1135; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_387;
  wire [388:0] _GEN_1136; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_388;
  wire [389:0] _GEN_1137; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_389;
  wire [390:0] _GEN_1138; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_390;
  wire [391:0] _GEN_1139; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_391;
  wire [392:0] _GEN_1140; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_392;
  wire [393:0] _GEN_1141; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_393;
  wire [394:0] _GEN_1142; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_394;
  wire [395:0] _GEN_1143; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_395;
  wire [396:0] _GEN_1144; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_396;
  wire [397:0] _GEN_1145; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_397;
  wire [398:0] _GEN_1146; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_398;
  wire [399:0] _GEN_1147; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_399;
  wire [400:0] _GEN_1148; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_400;
  wire [401:0] _GEN_1149; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_401;
  wire [402:0] _GEN_1150; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_402;
  wire [403:0] _GEN_1151; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_403;
  wire [404:0] _GEN_1152; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_404;
  wire [405:0] _GEN_1153; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_405;
  wire [406:0] _GEN_1154; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_406;
  wire [407:0] _GEN_1155; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_407;
  wire [408:0] _GEN_1156; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_408;
  wire [409:0] _GEN_1157; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_409;
  wire [410:0] _GEN_1158; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_410;
  wire [411:0] _GEN_1159; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_411;
  wire [412:0] _GEN_1160; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_412;
  wire [413:0] _GEN_1161; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_413;
  wire [414:0] _GEN_1162; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_414;
  wire [415:0] _GEN_1163; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_415;
  wire [416:0] _GEN_1164; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_416;
  wire [417:0] _GEN_1165; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_417;
  wire [418:0] _GEN_1166; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_418;
  wire [419:0] _GEN_1167; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_419;
  wire [420:0] _GEN_1168; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_420;
  wire [421:0] _GEN_1169; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_421;
  wire [422:0] _GEN_1170; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_422;
  wire [423:0] _GEN_1171; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_423;
  wire [424:0] _GEN_1172; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_424;
  wire [425:0] _GEN_1173; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_425;
  wire [426:0] _GEN_1174; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_426;
  wire [427:0] _GEN_1175; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_427;
  wire [428:0] _GEN_1176; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_428;
  wire [429:0] _GEN_1177; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_429;
  wire [430:0] _GEN_1178; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_430;
  wire [431:0] _GEN_1179; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_431;
  wire [432:0] _GEN_1180; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_432;
  wire [433:0] _GEN_1181; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_433;
  wire [434:0] _GEN_1182; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_434;
  wire [435:0] _GEN_1183; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_435;
  wire [436:0] _GEN_1184; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_436;
  wire [437:0] _GEN_1185; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_437;
  wire [438:0] _GEN_1186; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_438;
  wire [439:0] _GEN_1187; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_439;
  wire [440:0] _GEN_1188; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_440;
  wire [441:0] _GEN_1189; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_441;
  wire [442:0] _GEN_1190; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_442;
  wire [443:0] _GEN_1191; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_443;
  wire [444:0] _GEN_1192; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_444;
  wire [445:0] _GEN_1193; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_445;
  wire [446:0] _GEN_1194; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_446;
  wire [447:0] _GEN_1195; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_447;
  wire [448:0] _GEN_1196; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_448;
  wire [449:0] _GEN_1197; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_449;
  wire [450:0] _GEN_1198; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_450;
  wire [451:0] _GEN_1199; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_451;
  wire [452:0] _GEN_1200; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_452;
  wire [453:0] _GEN_1201; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_453;
  wire [454:0] _GEN_1202; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_454;
  wire [455:0] _GEN_1203; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_455;
  wire [456:0] _GEN_1204; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_456;
  wire [457:0] _GEN_1205; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_457;
  wire [458:0] _GEN_1206; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_458;
  wire [459:0] _GEN_1207; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_459;
  wire [460:0] _GEN_1208; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_460;
  wire [461:0] _GEN_1209; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_461;
  wire [462:0] _GEN_1210; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_462;
  wire [463:0] _GEN_1211; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_463;
  wire [464:0] _GEN_1212; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_464;
  wire [465:0] _GEN_1213; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_465;
  wire [466:0] _GEN_1214; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_466;
  wire [467:0] _GEN_1215; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_467;
  wire [468:0] _GEN_1216; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_468;
  wire [469:0] _GEN_1217; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_469;
  wire [470:0] _GEN_1218; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_470;
  wire [471:0] _GEN_1219; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_471;
  wire [472:0] _GEN_1220; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_472;
  wire [473:0] _GEN_1221; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_473;
  wire [474:0] _GEN_1222; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_474;
  wire [475:0] _GEN_1223; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_475;
  wire [476:0] _GEN_1224; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_476;
  wire [477:0] _GEN_1225; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_477;
  wire [478:0] _GEN_1226; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_478;
  wire [479:0] _GEN_1227; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_479;
  wire [480:0] _GEN_1228; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_480;
  wire [481:0] _GEN_1229; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_481;
  wire [482:0] _GEN_1230; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_482;
  wire [483:0] _GEN_1231; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_483;
  wire [484:0] _GEN_1232; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_484;
  wire [485:0] _GEN_1233; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_485;
  wire [486:0] _GEN_1234; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_486;
  wire [487:0] _GEN_1235; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_487;
  wire [488:0] _GEN_1236; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_488;
  wire [489:0] _GEN_1237; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_489;
  wire [490:0] _GEN_1238; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_490;
  wire [491:0] _GEN_1239; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_491;
  wire [492:0] _GEN_1240; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_492;
  wire [493:0] _GEN_1241; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_493;
  wire [494:0] _GEN_1242; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_494;
  wire [495:0] _GEN_1243; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_495;
  wire [496:0] _GEN_1244; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_496;
  wire [497:0] _GEN_1245; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_497;
  wire [498:0] _GEN_1246; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_498;
  wire [499:0] _GEN_1247; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_499;
  wire [500:0] _GEN_1248; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_500;
  wire [501:0] _GEN_1249; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_501;
  wire [502:0] _GEN_1250; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_502;
  wire [503:0] _GEN_1251; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_503;
  wire [504:0] _GEN_1252; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_504;
  wire [505:0] _GEN_1253; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_505;
  wire [506:0] _GEN_1254; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_506;
  wire [507:0] _GEN_1255; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_507;
  wire [508:0] _GEN_1256; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_508;
  wire [509:0] _GEN_1257; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_509;
  wire [510:0] _GEN_1258; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_510;
  wire [511:0] _GEN_1259; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_511;
  wire [512:0] _GEN_1260; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_512;
  wire [513:0] _GEN_1261; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_513;
  wire [514:0] _GEN_1262; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_514;
  wire [515:0] _GEN_1263; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_515;
  wire [516:0] _GEN_1264; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_516;
  wire [517:0] _GEN_1265; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_517;
  wire [518:0] _GEN_1266; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_518;
  wire [519:0] _GEN_1267; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_519;
  wire [520:0] _GEN_1268; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_520;
  wire [521:0] _GEN_1269; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_521;
  wire [522:0] _GEN_1270; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_522;
  wire [523:0] _GEN_1271; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_523;
  wire [524:0] _GEN_1272; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_524;
  wire [525:0] _GEN_1273; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_525;
  wire [526:0] _GEN_1274; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_526;
  wire [527:0] _GEN_1275; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_527;
  wire [528:0] _GEN_1276; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_528;
  wire [529:0] _GEN_1277; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_529;
  wire [530:0] _GEN_1278; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_530;
  wire [531:0] _GEN_1279; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_531;
  wire [532:0] _GEN_1280; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_532;
  wire [533:0] _GEN_1281; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_533;
  wire [534:0] _GEN_1282; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_534;
  wire [535:0] _GEN_1283; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_535;
  wire [536:0] _GEN_1284; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_536;
  wire [537:0] _GEN_1285; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_537;
  wire [538:0] _GEN_1286; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_538;
  wire [539:0] _GEN_1287; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_539;
  wire [540:0] _GEN_1288; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_540;
  wire [541:0] _GEN_1289; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_541;
  wire [542:0] _GEN_1290; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_542;
  wire [543:0] _GEN_1291; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_543;
  wire [544:0] _GEN_1292; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_544;
  wire [545:0] _GEN_1293; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_545;
  wire [546:0] _GEN_1294; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_546;
  wire [547:0] _GEN_1295; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_547;
  wire [548:0] _GEN_1296; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_548;
  wire [549:0] _GEN_1297; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_549;
  wire [550:0] _GEN_1298; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_550;
  wire [551:0] _GEN_1299; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_551;
  wire [552:0] _GEN_1300; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_552;
  wire [553:0] _GEN_1301; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_553;
  wire [554:0] _GEN_1302; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_554;
  wire [555:0] _GEN_1303; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_555;
  wire [556:0] _GEN_1304; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_556;
  wire [557:0] _GEN_1305; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_557;
  wire [558:0] _GEN_1306; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_558;
  wire [559:0] _GEN_1307; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_559;
  wire [560:0] _GEN_1308; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_560;
  wire [561:0] _GEN_1309; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_561;
  wire [562:0] _GEN_1310; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_562;
  wire [563:0] _GEN_1311; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_563;
  wire [564:0] _GEN_1312; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_564;
  wire [565:0] _GEN_1313; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_565;
  wire [566:0] _GEN_1314; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_566;
  wire [567:0] _GEN_1315; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_567;
  wire [568:0] _GEN_1316; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_568;
  wire [569:0] _GEN_1317; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_569;
  wire [570:0] _GEN_1318; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_570;
  wire [571:0] _GEN_1319; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_571;
  wire [572:0] _GEN_1320; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_572;
  wire [573:0] _GEN_1321; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_573;
  wire [574:0] _GEN_1322; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_574;
  wire [575:0] _GEN_1323; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_575;
  wire [576:0] _GEN_1324; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_576;
  wire [577:0] _GEN_1325; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_577;
  wire [578:0] _GEN_1326; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_578;
  wire [579:0] _GEN_1327; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_579;
  wire [580:0] _GEN_1328; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_580;
  wire [581:0] _GEN_1329; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_581;
  wire [582:0] _GEN_1330; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_582;
  wire [583:0] _GEN_1331; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_583;
  wire [584:0] _GEN_1332; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_584;
  wire [585:0] _GEN_1333; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_585;
  wire [586:0] _GEN_1334; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_586;
  wire [587:0] _GEN_1335; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_587;
  wire [588:0] _GEN_1336; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_588;
  wire [589:0] _GEN_1337; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_589;
  wire [590:0] _GEN_1338; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_590;
  wire [591:0] _GEN_1339; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_591;
  wire [592:0] _GEN_1340; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_592;
  wire [593:0] _GEN_1341; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_593;
  wire [594:0] _GEN_1342; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_594;
  wire [595:0] _GEN_1343; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_595;
  wire [596:0] _GEN_1344; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_596;
  wire [597:0] _GEN_1345; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_597;
  wire [598:0] _GEN_1346; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_598;
  wire [599:0] _GEN_1347; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_599;
  wire [600:0] _GEN_1348; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_600;
  wire [601:0] _GEN_1349; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_601;
  wire [602:0] _GEN_1350; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_602;
  wire [603:0] _GEN_1351; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_603;
  wire [604:0] _GEN_1352; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_604;
  wire [605:0] _GEN_1353; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_605;
  wire [606:0] _GEN_1354; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_606;
  wire [607:0] _GEN_1355; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_607;
  wire [608:0] _GEN_1356; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_608;
  wire [609:0] _GEN_1357; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_609;
  wire [610:0] _GEN_1358; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_610;
  wire [611:0] _GEN_1359; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_611;
  wire [612:0] _GEN_1360; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_612;
  wire [613:0] _GEN_1361; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_613;
  wire [614:0] _GEN_1362; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_614;
  wire [615:0] _GEN_1363; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_615;
  wire [616:0] _GEN_1364; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_616;
  wire [617:0] _GEN_1365; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_617;
  wire [618:0] _GEN_1366; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_618;
  wire [619:0] _GEN_1367; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_619;
  wire [620:0] _GEN_1368; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_620;
  wire [621:0] _GEN_1369; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_621;
  wire [622:0] _GEN_1370; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_622;
  wire [623:0] _GEN_1371; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_623;
  wire [624:0] _GEN_1372; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_624;
  wire [625:0] _GEN_1373; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_625;
  wire [626:0] _GEN_1374; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_626;
  wire [627:0] _GEN_1375; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_627;
  wire [628:0] _GEN_1376; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_628;
  wire [629:0] _GEN_1377; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_629;
  wire [630:0] _GEN_1378; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_630;
  wire [631:0] _GEN_1379; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_631;
  wire [632:0] _GEN_1380; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_632;
  wire [633:0] _GEN_1381; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_633;
  wire [634:0] _GEN_1382; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_634;
  wire [635:0] _GEN_1383; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_635;
  wire [636:0] _GEN_1384; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_636;
  wire [637:0] _GEN_1385; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_637;
  wire [638:0] _GEN_1386; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_638;
  wire [639:0] _GEN_1387; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_639;
  wire [640:0] _GEN_1388; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_640;
  wire [641:0] _GEN_1389; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_641;
  wire [642:0] _GEN_1390; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_642;
  wire [643:0] _GEN_1391; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_643;
  wire [644:0] _GEN_1392; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_644;
  wire [645:0] _GEN_1393; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_645;
  wire [646:0] _GEN_1394; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_646;
  wire [647:0] _GEN_1395; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_647;
  wire [648:0] _GEN_1396; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_648;
  wire [649:0] _GEN_1397; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_649;
  wire [650:0] _GEN_1398; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_650;
  wire [651:0] _GEN_1399; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_651;
  wire [652:0] _GEN_1400; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_652;
  wire [653:0] _GEN_1401; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_653;
  wire [654:0] _GEN_1402; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_654;
  wire [655:0] _GEN_1403; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_655;
  wire [656:0] _GEN_1404; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_656;
  wire [657:0] _GEN_1405; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_657;
  wire [658:0] _GEN_1406; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_658;
  wire [659:0] _GEN_1407; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_659;
  wire [660:0] _GEN_1408; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_660;
  wire [661:0] _GEN_1409; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_661;
  wire [662:0] _GEN_1410; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_662;
  wire [663:0] _GEN_1411; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_663;
  wire [664:0] _GEN_1412; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_664;
  wire [665:0] _GEN_1413; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_665;
  wire [666:0] _GEN_1414; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_666;
  wire [667:0] _GEN_1415; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_667;
  wire [668:0] _GEN_1416; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_668;
  wire [669:0] _GEN_1417; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_669;
  wire [670:0] _GEN_1418; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_670;
  wire [671:0] _GEN_1419; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_671;
  wire [672:0] _GEN_1420; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_672;
  wire [673:0] _GEN_1421; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_673;
  wire [674:0] _GEN_1422; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_674;
  wire [675:0] _GEN_1423; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_675;
  wire [676:0] _GEN_1424; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_676;
  wire [677:0] _GEN_1425; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_677;
  wire [678:0] _GEN_1426; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_678;
  wire [679:0] _GEN_1427; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_679;
  wire [680:0] _GEN_1428; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_680;
  wire [681:0] _GEN_1429; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_681;
  wire [682:0] _GEN_1430; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_682;
  wire [683:0] _GEN_1431; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_683;
  wire [684:0] _GEN_1432; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_684;
  wire [685:0] _GEN_1433; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_685;
  wire [686:0] _GEN_1434; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_686;
  wire [687:0] _GEN_1435; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_687;
  wire [688:0] _GEN_1436; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_688;
  wire [689:0] _GEN_1437; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_689;
  wire [690:0] _GEN_1438; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_690;
  wire [691:0] _GEN_1439; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_691;
  wire [692:0] _GEN_1440; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_692;
  wire [693:0] _GEN_1441; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_693;
  wire [694:0] _GEN_1442; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_694;
  wire [695:0] _GEN_1443; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_695;
  wire [696:0] _GEN_1444; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_696;
  wire [697:0] _GEN_1445; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_698;
  wire [698:0] _GEN_1446; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_699;
  wire [699:0] _GEN_1447; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_700;
  wire [700:0] _GEN_1448; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_701;
  wire [701:0] _GEN_1449; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_702;
  wire [702:0] _GEN_1450; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_703;
  wire [703:0] _GEN_1451; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_704;
  wire [704:0] _GEN_1452; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_705;
  wire [705:0] _GEN_1453; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_706;
  wire [706:0] _GEN_1454; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_707;
  wire [707:0] _GEN_1455; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_708;
  wire [708:0] _GEN_1456; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_709;
  wire [709:0] _GEN_1457; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_710;
  wire [710:0] _GEN_1458; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_711;
  wire [711:0] _GEN_1459; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_712;
  wire [712:0] _GEN_1460; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_713;
  wire [713:0] _GEN_1461; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_714;
  wire [714:0] _GEN_1462; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_715;
  wire [715:0] _GEN_1463; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_716;
  wire [716:0] _GEN_1464; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_717;
  wire [717:0] _GEN_1465; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_718;
  wire [718:0] _GEN_1466; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_719;
  wire [719:0] _GEN_1467; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_720;
  wire [720:0] _GEN_1468; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_721;
  wire [721:0] _GEN_1469; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_722;
  wire [722:0] _GEN_1470; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_723;
  wire [723:0] _GEN_1471; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_724;
  wire [724:0] _GEN_1472; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_725;
  wire [725:0] _GEN_1473; // @[:Sodor3Stage.fir@3963.2]
  wire [726:0] _GEN_1474; // @[:Sodor3Stage.fir@3963.2]
  wire [727:0] _GEN_1475; // @[:Sodor3Stage.fir@3963.2]
  wire [728:0] _GEN_1476; // @[:Sodor3Stage.fir@3963.2]
  wire [729:0] _GEN_1477; // @[:Sodor3Stage.fir@3963.2]
  wire [730:0] _GEN_1478; // @[:Sodor3Stage.fir@3963.2]
  wire [731:0] _GEN_1479; // @[:Sodor3Stage.fir@3963.2]
  wire [732:0] _GEN_1480; // @[:Sodor3Stage.fir@3963.2]
  wire [733:0] _GEN_1481; // @[:Sodor3Stage.fir@3963.2]
  wire [734:0] _GEN_1482; // @[:Sodor3Stage.fir@3963.2]
  wire [735:0] _GEN_1483; // @[:Sodor3Stage.fir@3963.2]
  wire [736:0] _GEN_1484; // @[:Sodor3Stage.fir@3963.2]
  wire [737:0] _GEN_1485; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_738;
  wire [738:0] _GEN_1486; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_739;
  wire [739:0] _GEN_1487; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_740;
  wire [740:0] _GEN_1488; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_741;
  wire [741:0] _GEN_1489; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_742;
  wire [742:0] _GEN_1490; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_743;
  wire [743:0] _GEN_1491; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_744;
  wire [744:0] _GEN_1492; // @[:Sodor3Stage.fir@3963.2]
  wire  profilePin_745;
  Core core ( // @[top.scala 26:26:Sodor3Stage.fir@3971.4]
    .metaReset(core_metaReset),
    .clock(core_clock),
    .reset(core_reset),
    .io_imem_req_bits_addr(core_io_imem_req_bits_addr),
    .io_imem_resp_bits_data(core_io_imem_resp_bits_data),
    .io_dmem_req_bits_addr(core_io_dmem_req_bits_addr),
    .io_dmem_req_bits_data(core_io_dmem_req_bits_data),
    .io_dmem_req_bits_fcn(core_io_dmem_req_bits_fcn),
    .io_dmem_req_bits_typ(core_io_dmem_req_bits_typ),
    .io_dmem_resp_bits_data(core_io_dmem_resp_bits_data),
    ._GEN_338(core__GEN_338),
    ._GEN_224(core__GEN_224),
    ._GEN_218(core__GEN_218),
    ._GEN_21(core__GEN_21),
    ._GEN_91(core__GEN_91),
    ._GEN_323(core__GEN_323),
    ._GEN_302(core__GEN_302),
    ._GEN_51(core__GEN_51),
    ._GEN_304(core__GEN_304),
    ._GEN_199(core__GEN_199),
    ._GEN_6(core__GEN_6),
    ._GEN_148(core__GEN_148),
    ._GEN_239(core__GEN_239),
    ._GEN_403(core__GEN_403),
    ._GEN_1(core__GEN_1),
    ._GEN_24(core__GEN_24),
    ._GEN_247(core__GEN_247),
    ._GEN_106(core__GEN_106),
    ._GEN_317(core__GEN_317),
    ._GEN_133(core__GEN_133),
    ._GEN_205(core__GEN_205),
    ._GEN_385(core__GEN_385),
    ._GEN_39(core__GEN_39),
    ._GEN_232(core__GEN_232),
    ._GEN_418(core__GEN_418),
    ._GEN_127(core__GEN_127),
    ._GEN_197(core__GEN_197),
    ._GEN_331(core__GEN_331),
    ._GEN_190(core__GEN_190),
    ._GEN_12(core__GEN_12),
    ._GEN_226(core__GEN_226),
    ._GEN_296(core__GEN_296),
    ._GEN_9_0(core__GEN_9_0),
    ._GEN_45(core__GEN_45),
    ._GEN_112(core__GEN_112),
    ._GEN_298(core__GEN_298),
    ._GEN_203(core__GEN_203),
    ._GEN_72(core__GEN_72),
    ._GEN_211(core__GEN_211),
    ._GEN_325(core__GEN_325),
    ._GEN_397(core__GEN_397),
    ._GEN_0(core__GEN_0),
    ._GEN_424(core__GEN_424),
    ._GEN_30(core__GEN_30),
    ._GEN_310(core__GEN_310),
    ._GEN_319(core__GEN_319),
    ._GEN_66(core__GEN_66),
    ._GEN_9_1(core__GEN_9_1),
    ._GEN_212(core__GEN_212),
    ._GEN_220(core__GEN_220),
    ._GEN_214(core__GEN_214),
    ._GEN_100(core__GEN_100),
    ._GEN_109(core__GEN_109),
    ._GEN_320(core__GEN_320),
    ._GEN_313(core__GEN_313),
    ._GEN_282(core__GEN_282),
    ._GEN_200(core__GEN_200),
    ._GEN_177(core__GEN_177),
    ._GEN_208(core__GEN_208),
    ._GEN_388(core__GEN_388),
    ._GEN_391(core__GEN_391),
    ._GEN_381(core__GEN_381),
    ._GEN_412(core__GEN_412),
    ._GEN_27(core__GEN_27),
    ._GEN_276(core__GEN_276),
    ._GEN_191(core__GEN_191),
    ._GEN_181(core__GEN_181),
    ._GEN_54(core__GEN_54),
    ._GEN_193(core__GEN_193),
    ._GEN_190_0(core__GEN_190_0),
    ._GEN_15(core__GEN_15),
    ._GEN_289(core__GEN_289),
    ._GEN_12_0(core__GEN_12_0),
    ._GEN_406(core__GEN_406),
    ._GEN_299(core__GEN_299),
    ._GEN_48(core__GEN_48),
    ._GEN_115(core__GEN_115),
    ._GEN_311(core__GEN_311),
    ._GEN_206(core__GEN_206),
    ._GEN_367(core__GEN_367),
    ._GEN_175(core__GEN_175),
    ._GEN_6_0(core__GEN_6_0),
    ._GEN_305(core__GEN_305),
    ._GEN_33(core__GEN_33),
    ._GEN_274(core__GEN_274),
    ._GEN_121(core__GEN_121),
    ._GEN_307(core__GEN_307),
    ._GEN_373(core__GEN_373),
    ._GEN_375(core__GEN_375),
    ._GEN_229(core__GEN_229),
    ._GEN_94(core__GEN_94),
    ._GEN_292(core__GEN_292),
    ._GEN_183(core__GEN_183),
    ._GEN_376(core__GEN_376),
    ._GEN_382(core__GEN_382),
    ._GEN_0_0(core__GEN_0_0),
    ._GEN_10(core__GEN_10),
    ._GEN_370(core__GEN_370),
    ._GEN_349(core__GEN_349),
    ._GEN_196(core__GEN_196),
    ._GEN_186(core__GEN_186),
    ._GEN_262(core__GEN_262),
    ._GEN_400(core__GEN_400),
    ._GEN_103(core__GEN_103),
    ._GEN_264(core__GEN_264),
    ._GEN_295(core__GEN_295),
    ._GEN_355(core__GEN_355),
    ._GEN_159(core__GEN_159),
    ._GEN_202(core__GEN_202),
    ._GEN_171(core__GEN_171),
    ._GEN_357(core__GEN_357),
    ._GEN_270(core__GEN_270),
    ._GEN_277(core__GEN_277),
    ._GEN_384(core__GEN_384),
    ._GEN_36(core__GEN_36),
    ._GEN_285(core__GEN_285),
    ._GEN_165(core__GEN_165),
    ._GEN_279(core__GEN_279),
    ._GEN_194(core__GEN_194),
    ._GEN_184(core__GEN_184),
    ._GEN_378(core__GEN_378),
    ._GEN_293(core__GEN_293),
    ._GEN_21_0(core__GEN_21_0),
    ._GEN_301(core__GEN_301),
    ._GEN_157(core__GEN_157),
    ._GEN_3_0(core__GEN_3_0),
    ._GEN_361(core__GEN_361),
    ._GEN_394(core__GEN_394),
    ._GEN_15_0(core__GEN_15_0),
    ._GEN_256(core__GEN_256),
    ._GEN_363(core__GEN_363),
    ._GEN_9_2(core__GEN_9_2),
    ._GEN_258(core__GEN_258),
    ._GEN_97(core__GEN_97),
    ._GEN_283(core__GEN_283),
    ._GEN_163(core__GEN_163),
    ._GEN_178(core__GEN_178),
    ._GEN_345(core__GEN_345),
    ._GEN_339(core__GEN_339),
    ._GEN_8(core__GEN_8),
    ._GEN_11(core__GEN_11),
    ._GEN_18(core__GEN_18),
    ._GEN_259(core__GEN_259),
    ._GEN_147(core__GEN_147),
    ._GEN_358(core__GEN_358),
    ._GEN_330(core__GEN_330),
    ._GEN_172(core__GEN_172),
    ._GEN_86(core__GEN_86),
    ._GEN_13(core__GEN_13),
    ._GEN_271(core__GEN_271),
    ._GEN_265(core__GEN_265),
    ._GEN_280(core__GEN_280),
    ._GEN_160(core__GEN_160),
    ._GEN_273(core__GEN_273),
    ._GEN_343(core__GEN_343),
    ._GEN_379(core__GEN_379),
    ._GEN_351(core__GEN_351),
    ._GEN_238(core__GEN_238),
    ._GEN_231(core__GEN_231),
    ._GEN_189(core__GEN_189),
    ._GEN_337(core__GEN_337),
    ._GEN_153(core__GEN_153),
    ._GEN_288(core__GEN_288),
    ._GEN_364(core__GEN_364),
    ._GEN_244(core__GEN_244),
    ._GEN_366(core__GEN_366),
    ._GEN_252(core__GEN_252),
    ._GEN_180(core__GEN_180),
    ._GEN_166(core__GEN_166),
    ._GEN_71(core__GEN_71),
    ._GEN_174(core__GEN_174),
    ._GEN_168(core__GEN_168),
    ._GEN_372(core__GEN_372),
    ._GEN_3_1(core__GEN_3_1),
    ._GEN_387(core__GEN_387),
    ._GEN_246(core__GEN_246),
    ._GEN_267(core__GEN_267),
    ._GEN_286(core__GEN_286),
    ._GEN_151(core__GEN_151),
    ._GEN_187(core__GEN_187),
    ._GEN_354(core__GEN_354),
    ._GEN_213(core__GEN_213),
    ._GEN_249(core__GEN_249),
    ._GEN_319_0(core__GEN_319_0),
    ._GEN_268(core__GEN_268),
    ._GEN_240(core__GEN_240),
    ._GEN_141(core__GEN_141),
    ._GEN_135(core__GEN_135),
    ._GEN_226_0(core__GEN_226_0),
    ._GEN_234(core__GEN_234),
    ._GEN_348(core__GEN_348),
    ._GEN_261(core__GEN_261),
    ._GEN_312(core__GEN_312),
    ._GEN_53(core__GEN_53),
    ._GEN_333(core__GEN_333),
    ._GEN_147_0(core__GEN_147_0),
    ._GEN_68(core__GEN_68),
    ._GEN_156(core__GEN_156),
    ._GEN_352(core__GEN_352),
    ._GEN_247_0(core__GEN_247_0),
    ._GEN_360(core__GEN_360),
    ._GEN_369(core__GEN_369),
    ._GEN_325_0(core__GEN_325_0),
    ._GEN_2(core__GEN_2),
    ._GEN_74(core__GEN_74),
    ._GEN_327(core__GEN_327),
    ._GEN_169(core__GEN_169),
    ._GEN_89(core__GEN_89),
    ._GEN_162(core__GEN_162),
    ._GEN_232_0(core__GEN_232_0),
    ._GEN_426(core__GEN_426),
    ._GEN_7_0(core__GEN_7_0),
    ._GEN_331_0(core__GEN_331_0),
    ._GEN_129(core__GEN_129),
    ._GEN_346(core__GEN_346),
    ._GEN_154(core__GEN_154),
    ._GEN_340(core__GEN_340),
    ._GEN_253(core__GEN_253),
    ._GEN_228(core__GEN_228),
    ._GEN_411(core__GEN_411),
    ._GEN_255(core__GEN_255),
    ._GEN_120(core__GEN_120),
    ._GEN_211_0(core__GEN_211_0),
    ._GEN_80(core__GEN_80),
    ._GEN_220_0(core__GEN_220_0),
    ._GEN_342(core__GEN_342),
    ._GEN_229_0(core__GEN_229_0),
    ._GEN_393(core__GEN_393),
    ._GEN_292_0(core__GEN_292_0),
    ._GEN_307_0(core__GEN_307_0),
    ._GEN_193_0(core__GEN_193_0),
    ._GEN_56(core__GEN_56),
    ._GEN_144(core__GEN_144),
    ._GEN_17(core__GEN_17),
    ._GEN_11_1(core__GEN_11_1),
    ._GEN_408(core__GEN_408),
    ._GEN_222(core__GEN_222),
    ._GEN_313_0(core__GEN_313_0),
    ._GEN_117(core__GEN_117),
    ._GEN_328(core__GEN_328),
    ._GEN_321(core__GEN_321),
    ._GEN_2_0(core__GEN_2_0),
    ._GEN_235(core__GEN_235),
    ._GEN_243(core__GEN_243),
    ._GEN_237(core__GEN_237),
    ._GEN_123(core__GEN_123),
    ._GEN_102(core__GEN_102),
    ._GEN_3_2(core__GEN_3_2),
    ._GEN_62(core__GEN_62),
    ._GEN_150(core__GEN_150),
    ._GEN_336(core__GEN_336),
    ._GEN_201(core__GEN_201),
    ._GEN_195(core__GEN_195),
    ._GEN_23(core__GEN_23),
    ._GEN_414(core__GEN_414),
    ._GEN_250(core__GEN_250),
    ._GEN_300(core__GEN_300),
    ._GEN_294(core__GEN_294),
    ._GEN_309(core__GEN_309),
    ._GEN_77(core__GEN_77),
    ._GEN_208_0(core__GEN_208_0),
    ._GEN_83(core__GEN_83),
    ._GEN_214_0(core__GEN_214_0),
    ._GEN_216(core__GEN_216),
    ._GEN_241(core__GEN_241),
    ._GEN_420(core__GEN_420),
    ._GEN_35(core__GEN_35),
    ._GEN_5_0(core__GEN_5_0),
    ._GEN_41(core__GEN_41),
    ._GEN_315(core__GEN_315),
    ._GEN_429(core__GEN_429),
    ._GEN_138(core__GEN_138),
    ._GEN_334(core__GEN_334),
    ._GEN_217(core__GEN_217),
    ._GEN_402(core__GEN_402),
    ._GEN_17_0(core__GEN_17_0),
    ._GEN_225(core__GEN_225),
    ._GEN_105(core__GEN_105),
    ._GEN_316(core__GEN_316),
    ._GEN_50(core__GEN_50),
    ._GEN_44(core__GEN_44),
    ._GEN_324(core__GEN_324),
    ._GEN_180_0(core__GEN_180_0),
    ._GEN_318(core__GEN_318),
    ._GEN_384_0(core__GEN_384_0),
    ._GEN_396(core__GEN_396),
    ._GEN_386(core__GEN_386),
    ._GEN_38(core__GEN_38),
    ._GEN_301_0(core__GEN_301_0),
    ._GEN_196_0(core__GEN_196_0),
    ._GEN_186_0(core__GEN_186_0),
    ._GEN_65(core__GEN_65),
    ._GEN_295_0(core__GEN_295_0),
    ._GEN_20(core__GEN_20),
    ._GEN_223(core__GEN_223),
    ._GEN_23_0(core__GEN_23_0),
    ._GEN_417(core__GEN_417),
    ._GEN_111(core__GEN_111),
    ._GEN_322(core__GEN_322),
    ._GEN_210(core__GEN_210),
    ._GEN_5_1(core__GEN_5_1),
    ._GEN_219(core__GEN_219),
    ._GEN_279_0(core__GEN_279_0),
    ._GEN_310_0(core__GEN_310_0),
    ._GEN_285_0(core__GEN_285_0),
    ._GEN_423(core__GEN_423),
    ._GEN_132(core__GEN_132),
    ._GEN_126(core__GEN_126),
    ._GEN_287(core__GEN_287),
    ._GEN_202_0(core__GEN_202_0),
    ._GEN_378_0(core__GEN_378_0),
    ._GEN_90(core__GEN_90),
    ._GEN_204(core__GEN_204),
    ._GEN_99(core__GEN_99),
    ._GEN_303(core__GEN_303),
    ._GEN_297(core__GEN_297),
    ._GEN_59(core__GEN_59),
    ._GEN_188(core__GEN_188),
    ._GEN_198(core__GEN_198),
    ._GEN_351_0(core__GEN_351_0),
    ._GEN_176(core__GEN_176),
    ._GEN_387_0(core__GEN_387_0),
    ._GEN_11_2(core__GEN_11_2),
    ._GEN_380(core__GEN_380),
    ._GEN_93(core__GEN_93),
    ._GEN_161(core__GEN_161),
    ._GEN_192(core__GEN_192),
    ._GEN_189_0(core__GEN_189_0),
    ._GEN_14_0(core__GEN_14_0),
    ._GEN_372_0(core__GEN_372_0),
    ._GEN_207(core__GEN_207),
    ._GEN_267_0(core__GEN_267_0),
    ._GEN_405(core__GEN_405),
    ._GEN_260(core__GEN_260),
    ._GEN_26(core__GEN_26),
    ._GEN_114(core__GEN_114),
    ._GEN_269(core__GEN_269),
    ._GEN_174_0(core__GEN_174_0),
    ._GEN_205_0(core__GEN_205_0),
    ._GEN_182(core__GEN_182),
    ._GEN_399(core__GEN_399),
    ._GEN_368(core__GEN_368),
    ._GEN_273_0(core__GEN_273_0),
    ._GEN_390(core__GEN_390),
    ._GEN_32(core__GEN_32),
    ._GEN_281(core__GEN_281),
    ._GEN_275(core__GEN_275),
    ._GEN_291(core__GEN_291),
    ._GEN_168_0(core__GEN_168_0),
    ._GEN_47(core__GEN_47),
    ._GEN_199_0(core__GEN_199_0),
    ._GEN_5_2(core__GEN_5_2),
    ._GEN_389(core__GEN_389),
    ._GEN_298_0(core__GEN_298_0),
    ._GEN_304_0(core__GEN_304_0),
    ._GEN_306(core__GEN_306),
    ._GEN_366_0(core__GEN_366_0),
    ._GEN_8_1(core__GEN_8_1),
    ._GEN_374(core__GEN_374),
    ._GEN_108(core__GEN_108),
    ._GEN_360_0(core__GEN_360_0),
    ._GEN_288_0(core__GEN_288_0),
    ._GEN_356(core__GEN_356),
    ._GEN_375_0(core__GEN_375_0),
    ._GEN_255_0(core__GEN_255_0),
    ._GEN_261_0(core__GEN_261_0),
    ._GEN_20_0(core__GEN_20_0),
    ._GEN_14_1(core__GEN_14_1),
    ._GEN_29(core__GEN_29),
    ._GEN_270_0(core__GEN_270_0),
    ._GEN_150_0(core__GEN_150_0),
    ._GEN_333_0(core__GEN_333_0),
    ._GEN_82(core__GEN_82),
    ._GEN_177_0(core__GEN_177_0),
    ._GEN_170(core__GEN_170),
    ._GEN_381_0(core__GEN_381_0),
    ._GEN_185(core__GEN_185),
    ._GEN_1_1(core__GEN_1_1),
    ._GEN_276_0(core__GEN_276_0),
    ._GEN_10_0(core__GEN_10_0),
    ._GEN_278(core__GEN_278),
    ._GEN_143(core__GEN_143),
    ._GEN_354_0(core__GEN_354_0),
    ._GEN_348_0(core__GEN_348_0),
    ._GEN_249_0(core__GEN_249_0),
    ._GEN_96(core__GEN_96),
    ._GEN_9_3(core__GEN_9_3),
    ._GEN_263(core__GEN_263),
    ._GEN_164(core__GEN_164),
    ._GEN_158(core__GEN_158),
    ._GEN_369_0(core__GEN_369_0),
    ._GEN_183_0(core__GEN_183_0),
    ._GEN_362(core__GEN_362),
    ._GEN_377(core__GEN_377),
    ._GEN_257(core__GEN_257),
    ._GEN_282_0(core__GEN_282_0),
    ._GEN_284(core__GEN_284),
    ._GEN_179(core__GEN_179),
    ._GEN_383(core__GEN_383),
    ._GEN_242(core__GEN_242),
    ._GEN_8_2(core__GEN_8_2),
    ._GEN_162_0(core__GEN_162_0),
    ._GEN_156_0(core__GEN_156_0),
    ._GEN_341(core__GEN_341),
    ._GEN_76(core__GEN_76),
    ._GEN_165_0(core__GEN_165_0),
    ._GEN_173(core__GEN_173),
    ._GEN_224_0(core__GEN_224_0),
    ._GEN_359(core__GEN_359),
    ._GEN_251(core__GEN_251),
    ._GEN_131(core__GEN_131),
    ._GEN_7_1(core__GEN_7_1),
    ._GEN_146(core__GEN_146),
    ._GEN_342_0(core__GEN_342_0),
    ._GEN_350(core__GEN_350),
    ._GEN_344(core__GEN_344),
    ._GEN_239_0(core__GEN_239_0),
    ._GEN_264_0(core__GEN_264_0),
    ._GEN_272(core__GEN_272),
    ._GEN_64(core__GEN_64),
    ._GEN_58(core__GEN_58),
    ._GEN_159_0(core__GEN_159_0),
    ._GEN_222_0(core__GEN_222_0),
    ._GEN_363_0(core__GEN_363_0),
    ._GEN_357_0(core__GEN_357_0),
    ._GEN_230(core__GEN_230),
    ._GEN_365(core__GEN_365),
    ._GEN_321_0(core__GEN_321_0),
    ._GEN_7_2(core__GEN_7_2),
    ._GEN_330_0(core__GEN_330_0),
    ._GEN_323_0(core__GEN_323_0),
    ._GEN_85(core__GEN_85),
    ._GEN_338_0(core__GEN_338_0),
    ._GEN_79(core__GEN_79),
    ._GEN_243_0(core__GEN_243_0),
    ._GEN_2_2(core__GEN_2_2),
    ._GEN_237_0(core__GEN_237_0),
    ._GEN_245(core__GEN_245),
    ._GEN_12_1(core__GEN_12_1),
    ._GEN_315_0(core__GEN_315_0),
    ._GEN_336_0(core__GEN_336_0),
    ._GEN_70(core__GEN_70),
    ._GEN_152(core__GEN_152),
    ._GEN_167(core__GEN_167),
    ._GEN_422(core__GEN_422),
    ._GEN_258_0(core__GEN_258_0),
    ._GEN_371(core__GEN_371),
    ._GEN_266(core__GEN_266),
    ._GEN_125(core__GEN_125),
    ._GEN_171_0(core__GEN_171_0),
    ._GEN_212_0(core__GEN_212_0),
    ._GEN_303_0(core__GEN_303_0),
    ._GEN_254(core__GEN_254),
    ._GEN_146_0(core__GEN_146_0),
    ._GEN_13_0(core__GEN_13_0),
    ._GEN_155(core__GEN_155),
    ._GEN_149(core__GEN_149),
    ._GEN_225_0(core__GEN_225_0),
    ._GEN_227(core__GEN_227),
    ._GEN_113(core__GEN_113),
    ._GEN_140(core__GEN_140),
    ._GEN_326(core__GEN_326),
    ._GEN_7_3(core__GEN_7_3),
    ._GEN_231_0(core__GEN_231_0),
    ._GEN_425(core__GEN_425),
    ._GEN_404(core__GEN_404),
    ._GEN_240_0(core__GEN_240_0),
    ._GEN_353(core__GEN_353),
    ._GEN_248(core__GEN_248),
    ._GEN_107(core__GEN_107),
    ._GEN_6_3(core__GEN_6_3),
    ._GEN_311_0(core__GEN_311_0),
    ._GEN_339_0(core__GEN_339_0),
    ._GEN_153_0(core__GEN_153_0),
    ._GEN_73(core__GEN_73),
    ._GEN_67(core__GEN_67),
    ._GEN_347(core__GEN_347),
    ._GEN_206_0(core__GEN_206_0),
    ._GEN_252_0(core__GEN_252_0),
    ._GEN_410(core__GEN_410),
    ._GEN_297_0(core__GEN_297_0),
    ._GEN_419(core__GEN_419),
    ._GEN_233(core__GEN_233),
    ._GEN_305_0(core__GEN_305_0),
    ._GEN_128(core__GEN_128),
    ._GEN_324_0(core__GEN_324_0),
    ._GEN_332(core__GEN_332),
    ._GEN_219_0(core__GEN_219_0),
    ._GEN_88(core__GEN_88),
    ._GEN_1_3(core__GEN_1_3),
    ._GEN_246_0(core__GEN_246_0),
    ._GEN_318_0(core__GEN_318_0),
    ._GEN_52(core__GEN_52),
    ._GEN_46(core__GEN_46),
    ._GEN_134(core__GEN_134),
    ._GEN_345_0(core__GEN_345_0),
    ._GEN_204_0(core__GEN_204_0),
    ._GEN_213_0(core__GEN_213_0),
    ._GEN_228_0(core__GEN_228_0),
    ._GEN_221(core__GEN_221),
    ._GEN_407(core__GEN_407),
    ._GEN_382_0(core__GEN_382_0),
    ._GEN_28(core__GEN_28),
    ._GEN_281_0(core__GEN_281_0),
    ._GEN_4_1(core__GEN_4_1),
    ._GEN_40(core__GEN_40),
    ._GEN_55(core__GEN_55),
    ._GEN_329(core__GEN_329),
    ._GEN_194_0(core__GEN_194_0),
    ._GEN_392(core__GEN_392),
    ._GEN_0_2(core__GEN_0_2),
    ._GEN_234_0(core__GEN_234_0),
    ._GEN_10_2(core__GEN_10_2),
    ._GEN_236(core__GEN_236),
    ._GEN_101(core__GEN_101),
    ._GEN_312_0(core__GEN_312_0),
    ._GEN_192_0(core__GEN_192_0),
    ._GEN_306_0(core__GEN_306_0),
    ._GEN_61(core__GEN_61),
    ._GEN_207_0(core__GEN_207_0),
    ._GEN_16(core__GEN_16),
    ._GEN_22(core__GEN_22),
    ._GEN_300_0(core__GEN_300_0),
    ._GEN_34(core__GEN_34),
    ._GEN_116(core__GEN_116),
    ._GEN_122(core__GEN_122),
    ._GEN_327_0(core__GEN_327_0),
    ._GEN_182_0(core__GEN_182_0),
    ._GEN_320_0(core__GEN_320_0),
    ._GEN_215(core__GEN_215),
    ._GEN_335(core__GEN_335),
    ._GEN_291_0(core__GEN_291_0),
    ._GEN_290(core__GEN_290),
    ._GEN_293_0(core__GEN_293_0),
    ._GEN_428(core__GEN_428),
    ._GEN_49(core__GEN_49),
    ._GEN_137(core__GEN_137),
    ._GEN_200_0(core__GEN_200_0),
    ._GEN_209(core__GEN_209),
    ._GEN_95(core__GEN_95),
    ._GEN_413(core__GEN_413),
    ._GEN_314(core__GEN_314),
    ._GEN_308(core__GEN_308),
    ._GEN_4_2(core__GEN_4_2),
    ._GEN_383_0(core__GEN_383_0),
    ._GEN_16_0(core__GEN_16_0),
    ._GEN_395(core__GEN_395),
    ._GEN_385_0(core__GEN_385_0),
    ._GEN_104(core__GEN_104),
    ._GEN_195_0(core__GEN_195_0),
    ._GEN_302_0(core__GEN_302_0),
    ._GEN_317_0(core__GEN_317_0),
    ._GEN_203_0(core__GEN_203_0),
    ._GEN_172_0(core__GEN_172_0),
    ._GEN_197_0(core__GEN_197_0),
    ._GEN_370_0(core__GEN_370_0),
    ._GEN_416(core__GEN_416),
    ._GEN_22_0(core__GEN_22_0),
    ._GEN_271_0(core__GEN_271_0),
    ._GEN_119(core__GEN_119),
    ._GEN_185_0(core__GEN_185_0),
    ._GEN_179_0(core__GEN_179_0),
    ._GEN_216_0(core__GEN_216_0),
    ._GEN_379_0(core__GEN_379_0),
    ._GEN_187_0(core__GEN_187_0),
    ._GEN_401(core__GEN_401),
    ._GEN_43(core__GEN_43),
    ._GEN_278_0(core__GEN_278_0),
    ._GEN_296_0(core__GEN_296_0),
    ._GEN_286_0(core__GEN_286_0),
    ._GEN_201_0(core__GEN_201_0),
    ._GEN_364_0(core__GEN_364_0),
    ._GEN_1_4(core__GEN_1_4),
    ._GEN_210_0(core__GEN_210_0),
    ._GEN_98(core__GEN_98),
    ._GEN_263_0(core__GEN_263_0),
    ._GEN_309_0(core__GEN_309_0),
    ._GEN_37(core__GEN_37),
    ._GEN_164_0(core__GEN_164_0),
    ._GEN_110(core__GEN_110),
    ._GEN_362_0(core__GEN_362_0),
    ._GEN_19(core__GEN_19),
    ._GEN_377_0(core__GEN_377_0),
    ._GEN_218_0(core__GEN_218_0),
    ._GEN_294_0(core__GEN_294_0),
    ._GEN_284_0(core__GEN_284_0),
    ._GEN_371_0(core__GEN_371_0),
    ._GEN_260_0(core__GEN_260_0),
    ._GEN_266_0(core__GEN_266_0),
    ._GEN_380_0(core__GEN_380_0),
    ._GEN_25(core__GEN_25),
    ._GEN_365_0(core__GEN_365_0),
    ._GEN_181_0(core__GEN_181_0),
    ._GEN_175_0(core__GEN_175_0),
    ._GEN_251_0(core__GEN_251_0),
    ._GEN_15_1(core__GEN_15_1),
    ._GEN_289_0(core__GEN_289_0),
    ._GEN_359_0(core__GEN_359_0),
    ._GEN_352_0(core__GEN_352_0),
    ._GEN_14_2(core__GEN_14_2),
    ._GEN_152_0(core__GEN_152_0),
    ._GEN_31(core__GEN_31),
    ._GEN_274_0(core__GEN_274_0),
    ._GEN_160_0(core__GEN_160_0),
    ._GEN_169_0(core__GEN_169_0),
    ._GEN_191_0(core__GEN_191_0),
    ._GEN_188_0(core__GEN_188_0),
    ._GEN_373_0(core__GEN_373_0),
    ._GEN_19_0(core__GEN_19_0),
    ._GEN_367_0(core__GEN_367_0),
    ._GEN_268_0(core__GEN_268_0),
    ._GEN_173_0(core__GEN_173_0),
    ._GEN_290_0(core__GEN_290_0),
    ._GEN_280_0(core__GEN_280_0),
    ._GEN_287_0(core__GEN_287_0),
    ._GEN_154_0(core__GEN_154_0),
    ._GEN_87(core__GEN_87),
    ._GEN_299_0(core__GEN_299_0),
    ._GEN_386_0(core__GEN_386_0),
    ._GEN_10_3(core__GEN_10_3),
    ._GEN_245_0(core__GEN_245_0),
    ._GEN_398(core__GEN_398),
    ._GEN_4_3(core__GEN_4_3),
    ._GEN_388_0(core__GEN_388_0),
    ._GEN_253_0(core__GEN_253_0),
    ._GEN_92(core__GEN_92),
    ._GEN_5_3(core__GEN_5_3),
    ._GEN_272_0(core__GEN_272_0),
    ._GEN_344_0(core__GEN_344_0),
    ._GEN_198_0(core__GEN_198_0),
    ._GEN_167_0(core__GEN_167_0),
    ._GEN_346_0(core__GEN_346_0),
    ._GEN_334_0(core__GEN_334_0),
    ._GEN_340_0(core__GEN_340_0),
    ._GEN_254_0(core__GEN_254_0),
    ._GEN_13_2(core__GEN_13_2),
    ._GEN_3_4(core__GEN_3_4),
    ._GEN_256_0(core__GEN_256_0),
    ._GEN_328_0(core__GEN_328_0),
    ._GEN_161_0(core__GEN_161_0),
    ._GEN_347_0(core__GEN_347_0),
    ._GEN_81(core__GEN_81),
    ._GEN_355_0(core__GEN_355_0),
    ._GEN_170_0(core__GEN_170_0),
    ._GEN_7_5(core__GEN_7_5),
    ._GEN_8_3(core__GEN_8_3),
    ._GEN_275_0(core__GEN_275_0),
    ._GEN_269_0(core__GEN_269_0),
    ._GEN_155_0(core__GEN_155_0),
    ._GEN_277_0(core__GEN_277_0),
    ._GEN_69(core__GEN_69),
    ._GEN_157_0(core__GEN_157_0),
    ._GEN_368_0(core__GEN_368_0),
    ._GEN_233_0(core__GEN_233_0),
    ._GEN_227_0(core__GEN_227_0),
    ._GEN_235_0(core__GEN_235_0),
    ._GEN_184_0(core__GEN_184_0),
    ._GEN_326_0(core__GEN_326_0),
    ._GEN_149_0(core__GEN_149_0),
    ._GEN_60(core__GEN_60),
    ._GEN_283_0(core__GEN_283_0),
    ._GEN_142(core__GEN_142),
    ._GEN_353_0(core__GEN_353_0),
    ._GEN_178_0(core__GEN_178_0),
    ._GEN_248_0(core__GEN_248_0),
    ._GEN_241_0(core__GEN_241_0),
    ._GEN_361_0(core__GEN_361_0),
    ._GEN_136(core__GEN_136),
    ._GEN_75(core__GEN_75),
    ._GEN_163_0(core__GEN_163_0),
    ._GEN_349_0(core__GEN_349_0),
    ._GEN_374_0(core__GEN_374_0),
    ._GEN_427(core__GEN_427),
    ._GEN_376_0(core__GEN_376_0),
    ._GEN_262_0(core__GEN_262_0),
    ._GEN_332_0(core__GEN_332_0),
    ._GEN_176_0(core__GEN_176_0),
    ._GEN_166_0(core__GEN_166_0),
    ._GEN_358_0(core__GEN_358_0),
    ._GEN_314_0(core__GEN_314_0),
    ._GEN_308_0(core__GEN_308_0),
    ._GEN_42(core__GEN_42),
    ._GEN_265_0(core__GEN_265_0),
    ._GEN_316_0(core__GEN_316_0),
    ._GEN_130(core__GEN_130),
    ._GEN_124(core__GEN_124),
    ._GEN_341_0(core__GEN_341_0),
    ._GEN_343_0(core__GEN_343_0),
    ._GEN_223_0(core__GEN_223_0),
    ._GEN_238_0(core__GEN_238_0),
    ._GEN_118(core__GEN_118),
    ._GEN_5_4(core__GEN_5_4),
    ._GEN_151_0(core__GEN_151_0),
    ._GEN_145(core__GEN_145),
    ._GEN_337_0(core__GEN_337_0),
    ._GEN_18_0(core__GEN_18_0),
    ._GEN_356_0(core__GEN_356_0),
    ._GEN_244_0(core__GEN_244_0),
    ._GEN_409(core__GEN_409),
    ._GEN_11_3(core__GEN_11_3),
    ._GEN_322_0(core__GEN_322_0),
    ._GEN_158_0(core__GEN_158_0),
    ._GEN_209_0(core__GEN_209_0),
    ._GEN_78(core__GEN_78),
    ._GEN_217_0(core__GEN_217_0),
    ._GEN_221_0(core__GEN_221_0),
    ._GEN_236_0(core__GEN_236_0),
    ._GEN_421(core__GEN_421),
    ._GEN_415(core__GEN_415),
    ._GEN_335_0(core__GEN_335_0),
    ._GEN_329_0(core__GEN_329_0),
    ._GEN_63(core__GEN_63),
    ._GEN_230_0(core__GEN_230_0),
    ._GEN_242_0(core__GEN_242_0),
    ._GEN_257_0(core__GEN_257_0),
    ._GEN_6_4(core__GEN_6_4),
    ._GEN_57(core__GEN_57),
    ._GEN_250_0(core__GEN_250_0),
    ._GEN_259_0(core__GEN_259_0),
    ._GEN_139(core__GEN_139),
    ._GEN_350_0(core__GEN_350_0),
    ._GEN_215_0(core__GEN_215_0),
    ._GEN_84(core__GEN_84)
  );
  SyncScratchPadMemory memory ( // @[top.scala 29:28:Sodor3Stage.fir@3974.4]
    .metaReset(memory_metaReset),
    .clock(memory_clock),
    .io_core_ports_0_req_bits_addr(memory_io_core_ports_0_req_bits_addr),
    .io_core_ports_0_req_bits_data(memory_io_core_ports_0_req_bits_data),
    .io_core_ports_0_req_bits_fcn(memory_io_core_ports_0_req_bits_fcn),
    .io_core_ports_0_req_bits_typ(memory_io_core_ports_0_req_bits_typ),
    .io_core_ports_0_resp_bits_data(memory_io_core_ports_0_resp_bits_data),
    ._GEN_3_0(memory__GEN_3_0),
    ._GEN_7_0(memory__GEN_7_0),
    ._GEN_1_1(memory__GEN_1_1),
    ._GEN_4_0(memory__GEN_4_0),
    ._GEN_2_2(memory__GEN_2_2),
    ._GEN_3_4(memory__GEN_3_4),
    ._GEN_6_3(memory__GEN_6_3),
    ._GEN_0_2(memory__GEN_0_2),
    ._GEN_1_3(memory__GEN_1_3),
    ._GEN_2_4(memory__GEN_2_4),
    ._GEN_0_4(memory__GEN_0_4),
    ._GEN_5_6(memory__GEN_5_6)
  );
  assign core_metaReset = metaReset;
  assign memory_metaReset = metaReset;
  assign profilePin = core__GEN_1;
  assign profilePin_0 = core__GEN_5_3;
  assign _GEN_749 = {profilePin,profilePin_0}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_1 = core__GEN_6_3;
  assign _GEN_750 = {_GEN_749,profilePin_1}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_2 = core__GEN_7_0;
  assign _GEN_751 = {_GEN_750,profilePin_2}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_3 = core__GEN_8_3;
  assign _GEN_752 = {_GEN_751,profilePin_3}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_4 = core__GEN_9_3;
  assign _GEN_753 = {_GEN_752,profilePin_4}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_5 = core__GEN_10;
  assign _GEN_754 = {_GEN_753,profilePin_5}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_6 = core__GEN_11_3;
  assign _GEN_755 = {_GEN_754,profilePin_6}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_7 = core__GEN_12_1;
  assign _GEN_756 = {_GEN_755,profilePin_7}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_8 = core__GEN_13;
  assign _GEN_757 = {_GEN_756,profilePin_8}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_9 = core__GEN_14_2;
  assign _GEN_758 = {_GEN_757,profilePin_9}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_10 = core__GEN_0_0;
  assign _GEN_759 = {_GEN_758,profilePin_10}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_11 = core__GEN_1_4;
  assign _GEN_760 = {_GEN_759,profilePin_11}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_12 = core__GEN_2_2;
  assign _GEN_761 = {_GEN_760,profilePin_12}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_13 = core__GEN_3_1;
  assign _GEN_762 = {_GEN_761,profilePin_13}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_14 = core__GEN_4_3;
  assign _GEN_763 = {_GEN_762,profilePin_14}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_15 = core__GEN_5_2;
  assign _GEN_764 = {_GEN_763,profilePin_15}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_16 = core__GEN_6_0;
  assign _GEN_765 = {_GEN_764,profilePin_16}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_17 = core__GEN_7_5;
  assign _GEN_766 = {_GEN_765,profilePin_17}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_18 = core__GEN_8_2;
  assign _GEN_767 = {_GEN_766,profilePin_18}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_19 = core__GEN_9_2;
  assign _GEN_768 = {_GEN_767,profilePin_19}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_20 = core__GEN_10_3;
  assign _GEN_769 = {_GEN_768,profilePin_20}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_21 = core__GEN_11_2;
  assign _GEN_770 = {_GEN_769,profilePin_21}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_22 = core__GEN_12_0;
  assign _GEN_771 = {_GEN_770,profilePin_22}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_23 = core__GEN_13_2;
  assign _GEN_772 = {_GEN_771,profilePin_23}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_24 = core__GEN_14_1;
  assign _GEN_773 = {_GEN_772,profilePin_24}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_25 = core__GEN_15_0;
  assign _GEN_774 = {_GEN_773,profilePin_25}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_26 = core__GEN_16_0;
  assign _GEN_775 = {_GEN_774,profilePin_26}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_27 = core__GEN_17_0;
  assign _GEN_776 = {_GEN_775,profilePin_27}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_28 = core__GEN_18;
  assign _GEN_777 = {_GEN_776,profilePin_28}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_29 = core__GEN_19_0;
  assign _GEN_778 = {_GEN_777,profilePin_29}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_30 = core__GEN_20_0;
  assign _GEN_779 = {_GEN_778,profilePin_30}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_31 = core__GEN_21_0;
  assign _GEN_780 = {_GEN_779,profilePin_31}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_32 = core__GEN_22_0;
  assign _GEN_781 = {_GEN_780,profilePin_32}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_33 = core__GEN_23_0;
  assign _GEN_782 = {_GEN_781,profilePin_33}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_34 = core__GEN_24;
  assign _GEN_783 = {_GEN_782,profilePin_34}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_35 = core__GEN_25;
  assign _GEN_784 = {_GEN_783,profilePin_35}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_36 = core__GEN_26;
  assign _GEN_785 = {_GEN_784,profilePin_36}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_37 = core__GEN_27;
  assign _GEN_786 = {_GEN_785,profilePin_37}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_38 = core__GEN_28;
  assign _GEN_787 = {_GEN_786,profilePin_38}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_39 = core__GEN_29;
  assign _GEN_788 = {_GEN_787,profilePin_39}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_40 = core__GEN_30;
  assign _GEN_789 = {_GEN_788,profilePin_40}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_41 = core__GEN_31;
  assign _GEN_790 = {_GEN_789,profilePin_41}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_42 = core__GEN_32;
  assign _GEN_791 = {_GEN_790,profilePin_42}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_43 = core__GEN_33;
  assign _GEN_792 = {_GEN_791,profilePin_43}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_44 = core__GEN_34;
  assign _GEN_793 = {_GEN_792,profilePin_44}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_45 = core__GEN_35;
  assign _GEN_794 = {_GEN_793,profilePin_45}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_46 = core__GEN_36;
  assign _GEN_795 = {_GEN_794,profilePin_46}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_47 = core__GEN_37;
  assign _GEN_796 = {_GEN_795,profilePin_47}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_48 = core__GEN_38;
  assign _GEN_797 = {_GEN_796,profilePin_48}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_49 = core__GEN_39;
  assign _GEN_798 = {_GEN_797,profilePin_49}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_50 = core__GEN_40;
  assign _GEN_799 = {_GEN_798,profilePin_50}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_51 = core__GEN_41;
  assign _GEN_800 = {_GEN_799,profilePin_51}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_52 = core__GEN_42;
  assign _GEN_801 = {_GEN_800,profilePin_52}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_53 = core__GEN_43;
  assign _GEN_802 = {_GEN_801,profilePin_53}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_54 = core__GEN_44;
  assign _GEN_803 = {_GEN_802,profilePin_54}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_55 = core__GEN_45;
  assign _GEN_804 = {_GEN_803,profilePin_55}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_56 = core__GEN_46;
  assign _GEN_805 = {_GEN_804,profilePin_56}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_57 = core__GEN_47;
  assign _GEN_806 = {_GEN_805,profilePin_57}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_58 = core__GEN_48;
  assign _GEN_807 = {_GEN_806,profilePin_58}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_59 = core__GEN_49;
  assign _GEN_808 = {_GEN_807,profilePin_59}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_60 = core__GEN_50;
  assign _GEN_809 = {_GEN_808,profilePin_60}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_61 = core__GEN_51;
  assign _GEN_810 = {_GEN_809,profilePin_61}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_62 = core__GEN_52;
  assign _GEN_811 = {_GEN_810,profilePin_62}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_63 = core__GEN_53;
  assign _GEN_812 = {_GEN_811,profilePin_63}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_64 = core__GEN_54;
  assign _GEN_813 = {_GEN_812,profilePin_64}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_65 = core__GEN_55;
  assign _GEN_814 = {_GEN_813,profilePin_65}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_66 = core__GEN_56;
  assign _GEN_815 = {_GEN_814,profilePin_66}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_67 = core__GEN_57;
  assign _GEN_816 = {_GEN_815,profilePin_67}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_68 = core__GEN_58;
  assign _GEN_817 = {_GEN_816,profilePin_68}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_69 = core__GEN_59;
  assign _GEN_818 = {_GEN_817,profilePin_69}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_70 = core__GEN_60;
  assign _GEN_819 = {_GEN_818,profilePin_70}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_71 = core__GEN_61;
  assign _GEN_820 = {_GEN_819,profilePin_71}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_72 = core__GEN_62;
  assign _GEN_821 = {_GEN_820,profilePin_72}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_73 = core__GEN_63;
  assign _GEN_822 = {_GEN_821,profilePin_73}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_74 = core__GEN_64;
  assign _GEN_823 = {_GEN_822,profilePin_74}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_75 = core__GEN_65;
  assign _GEN_824 = {_GEN_823,profilePin_75}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_76 = core__GEN_66;
  assign _GEN_825 = {_GEN_824,profilePin_76}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_77 = core__GEN_67;
  assign _GEN_826 = {_GEN_825,profilePin_77}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_78 = core__GEN_68;
  assign _GEN_827 = {_GEN_826,profilePin_78}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_79 = core__GEN_69;
  assign _GEN_828 = {_GEN_827,profilePin_79}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_80 = core__GEN_70;
  assign _GEN_829 = {_GEN_828,profilePin_80}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_81 = core__GEN_71;
  assign _GEN_830 = {_GEN_829,profilePin_81}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_82 = core__GEN_72;
  assign _GEN_831 = {_GEN_830,profilePin_82}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_83 = core__GEN_73;
  assign _GEN_832 = {_GEN_831,profilePin_83}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_84 = core__GEN_74;
  assign _GEN_833 = {_GEN_832,profilePin_84}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_85 = core__GEN_75;
  assign _GEN_834 = {_GEN_833,profilePin_85}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_86 = core__GEN_76;
  assign _GEN_835 = {_GEN_834,profilePin_86}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_87 = core__GEN_77;
  assign _GEN_836 = {_GEN_835,profilePin_87}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_88 = core__GEN_78;
  assign _GEN_837 = {_GEN_836,profilePin_88}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_89 = core__GEN_79;
  assign _GEN_838 = {_GEN_837,profilePin_89}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_90 = core__GEN_80;
  assign _GEN_839 = {_GEN_838,profilePin_90}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_91 = core__GEN_81;
  assign _GEN_840 = {_GEN_839,profilePin_91}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_92 = core__GEN_82;
  assign _GEN_841 = {_GEN_840,profilePin_92}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_93 = core__GEN_83;
  assign _GEN_842 = {_GEN_841,profilePin_93}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_94 = core__GEN_84;
  assign _GEN_843 = {_GEN_842,profilePin_94}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_95 = core__GEN_85;
  assign _GEN_844 = {_GEN_843,profilePin_95}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_96 = core__GEN_86;
  assign _GEN_845 = {_GEN_844,profilePin_96}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_97 = core__GEN_87;
  assign _GEN_846 = {_GEN_845,profilePin_97}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_98 = core__GEN_88;
  assign _GEN_847 = {_GEN_846,profilePin_98}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_99 = core__GEN_89;
  assign _GEN_848 = {_GEN_847,profilePin_99}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_100 = core__GEN_90;
  assign _GEN_849 = {_GEN_848,profilePin_100}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_101 = core__GEN_91;
  assign _GEN_850 = {_GEN_849,profilePin_101}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_102 = core__GEN_92;
  assign _GEN_851 = {_GEN_850,profilePin_102}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_103 = core__GEN_93;
  assign _GEN_852 = {_GEN_851,profilePin_103}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_104 = core__GEN_94;
  assign _GEN_853 = {_GEN_852,profilePin_104}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_105 = core__GEN_95;
  assign _GEN_854 = {_GEN_853,profilePin_105}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_106 = core__GEN_96;
  assign _GEN_855 = {_GEN_854,profilePin_106}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_107 = core__GEN_97;
  assign _GEN_856 = {_GEN_855,profilePin_107}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_108 = core__GEN_98;
  assign _GEN_857 = {_GEN_856,profilePin_108}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_109 = core__GEN_99;
  assign _GEN_858 = {_GEN_857,profilePin_109}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_110 = core__GEN_100;
  assign _GEN_859 = {_GEN_858,profilePin_110}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_111 = core__GEN_101;
  assign _GEN_860 = {_GEN_859,profilePin_111}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_112 = core__GEN_102;
  assign _GEN_861 = {_GEN_860,profilePin_112}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_113 = core__GEN_103;
  assign _GEN_862 = {_GEN_861,profilePin_113}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_114 = core__GEN_104;
  assign _GEN_863 = {_GEN_862,profilePin_114}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_115 = core__GEN_105;
  assign _GEN_864 = {_GEN_863,profilePin_115}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_116 = core__GEN_106;
  assign _GEN_865 = {_GEN_864,profilePin_116}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_117 = core__GEN_107;
  assign _GEN_866 = {_GEN_865,profilePin_117}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_118 = core__GEN_108;
  assign _GEN_867 = {_GEN_866,profilePin_118}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_119 = core__GEN_109;
  assign _GEN_868 = {_GEN_867,profilePin_119}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_120 = core__GEN_110;
  assign _GEN_869 = {_GEN_868,profilePin_120}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_121 = core__GEN_111;
  assign _GEN_870 = {_GEN_869,profilePin_121}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_122 = core__GEN_112;
  assign _GEN_871 = {_GEN_870,profilePin_122}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_123 = core__GEN_113;
  assign _GEN_872 = {_GEN_871,profilePin_123}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_124 = core__GEN_114;
  assign _GEN_873 = {_GEN_872,profilePin_124}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_125 = core__GEN_115;
  assign _GEN_874 = {_GEN_873,profilePin_125}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_126 = core__GEN_116;
  assign _GEN_875 = {_GEN_874,profilePin_126}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_127 = core__GEN_117;
  assign _GEN_876 = {_GEN_875,profilePin_127}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_128 = core__GEN_118;
  assign _GEN_877 = {_GEN_876,profilePin_128}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_129 = core__GEN_119;
  assign _GEN_878 = {_GEN_877,profilePin_129}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_130 = core__GEN_120;
  assign _GEN_879 = {_GEN_878,profilePin_130}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_131 = core__GEN_121;
  assign _GEN_880 = {_GEN_879,profilePin_131}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_132 = core__GEN_122;
  assign _GEN_881 = {_GEN_880,profilePin_132}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_133 = core__GEN_123;
  assign _GEN_882 = {_GEN_881,profilePin_133}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_134 = core__GEN_124;
  assign _GEN_883 = {_GEN_882,profilePin_134}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_135 = core__GEN_125;
  assign _GEN_884 = {_GEN_883,profilePin_135}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_136 = core__GEN_126;
  assign _GEN_885 = {_GEN_884,profilePin_136}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_137 = core__GEN_127;
  assign _GEN_886 = {_GEN_885,profilePin_137}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_138 = core__GEN_128;
  assign _GEN_887 = {_GEN_886,profilePin_138}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_139 = core__GEN_129;
  assign _GEN_888 = {_GEN_887,profilePin_139}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_140 = core__GEN_130;
  assign _GEN_889 = {_GEN_888,profilePin_140}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_141 = core__GEN_131;
  assign _GEN_890 = {_GEN_889,profilePin_141}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_142 = core__GEN_132;
  assign _GEN_891 = {_GEN_890,profilePin_142}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_143 = core__GEN_133;
  assign _GEN_892 = {_GEN_891,profilePin_143}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_144 = core__GEN_134;
  assign _GEN_893 = {_GEN_892,profilePin_144}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_145 = core__GEN_135;
  assign _GEN_894 = {_GEN_893,profilePin_145}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_146 = core__GEN_136;
  assign _GEN_895 = {_GEN_894,profilePin_146}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_147 = core__GEN_137;
  assign _GEN_896 = {_GEN_895,profilePin_147}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_148 = core__GEN_138;
  assign _GEN_897 = {_GEN_896,profilePin_148}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_149 = core__GEN_139;
  assign _GEN_898 = {_GEN_897,profilePin_149}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_150 = core__GEN_140;
  assign _GEN_899 = {_GEN_898,profilePin_150}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_151 = core__GEN_141;
  assign _GEN_900 = {_GEN_899,profilePin_151}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_152 = core__GEN_142;
  assign _GEN_901 = {_GEN_900,profilePin_152}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_153 = core__GEN_143;
  assign _GEN_902 = {_GEN_901,profilePin_153}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_154 = core__GEN_144;
  assign _GEN_903 = {_GEN_902,profilePin_154}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_155 = core__GEN_145;
  assign _GEN_904 = {_GEN_903,profilePin_155}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_156 = core__GEN_146;
  assign _GEN_905 = {_GEN_904,profilePin_156}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_157 = core__GEN_147;
  assign _GEN_906 = {_GEN_905,profilePin_157}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_158 = core__GEN_148;
  assign _GEN_907 = {_GEN_906,profilePin_158}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_159 = core__GEN_149;
  assign _GEN_908 = {_GEN_907,profilePin_159}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_160 = core__GEN_150;
  assign _GEN_909 = {_GEN_908,profilePin_160}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_161 = core__GEN_151_0;
  assign _GEN_910 = {_GEN_909,profilePin_161}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_162 = core__GEN_152;
  assign _GEN_911 = {_GEN_910,profilePin_162}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_163 = core__GEN_153;
  assign _GEN_912 = {_GEN_911,profilePin_163}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_164 = core__GEN_154_0;
  assign _GEN_913 = {_GEN_912,profilePin_164}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_165 = core__GEN_155;
  assign _GEN_914 = {_GEN_913,profilePin_165}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_166 = core__GEN_156;
  assign _GEN_915 = {_GEN_914,profilePin_166}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_167 = core__GEN_157_0;
  assign _GEN_916 = {_GEN_915,profilePin_167}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_168 = core__GEN_158;
  assign _GEN_917 = {_GEN_916,profilePin_168}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_169 = core__GEN_159;
  assign _GEN_918 = {_GEN_917,profilePin_169}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_170 = core__GEN_160_0;
  assign _GEN_919 = {_GEN_918,profilePin_170}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_171 = core__GEN_161;
  assign _GEN_920 = {_GEN_919,profilePin_171}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_172 = core__GEN_162;
  assign _GEN_921 = {_GEN_920,profilePin_172}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_173 = core__GEN_163_0;
  assign _GEN_922 = {_GEN_921,profilePin_173}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_174 = core__GEN_164;
  assign _GEN_923 = {_GEN_922,profilePin_174}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_175 = core__GEN_165;
  assign _GEN_924 = {_GEN_923,profilePin_175}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_176 = core__GEN_166_0;
  assign _GEN_925 = {_GEN_924,profilePin_176}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_177 = core__GEN_167;
  assign _GEN_926 = {_GEN_925,profilePin_177}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_178 = core__GEN_168;
  assign _GEN_927 = {_GEN_926,profilePin_178}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_179 = core__GEN_169_0;
  assign _GEN_928 = {_GEN_927,profilePin_179}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_180 = core__GEN_170;
  assign _GEN_929 = {_GEN_928,profilePin_180}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_181 = core__GEN_171;
  assign _GEN_930 = {_GEN_929,profilePin_181}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_182 = core__GEN_172_0;
  assign _GEN_931 = {_GEN_930,profilePin_182}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_183 = core__GEN_173;
  assign _GEN_932 = {_GEN_931,profilePin_183}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_184 = core__GEN_174;
  assign _GEN_933 = {_GEN_932,profilePin_184}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_185 = core__GEN_175_0;
  assign _GEN_934 = {_GEN_933,profilePin_185}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_186 = core__GEN_176;
  assign _GEN_935 = {_GEN_934,profilePin_186}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_187 = core__GEN_177;
  assign _GEN_936 = {_GEN_935,profilePin_187}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_188 = core__GEN_178_0;
  assign _GEN_937 = {_GEN_936,profilePin_188}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_189 = core__GEN_179;
  assign _GEN_938 = {_GEN_937,profilePin_189}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_190 = core__GEN_180;
  assign _GEN_939 = {_GEN_938,profilePin_190}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_191 = core__GEN_181_0;
  assign _GEN_940 = {_GEN_939,profilePin_191}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_192 = core__GEN_182;
  assign _GEN_941 = {_GEN_940,profilePin_192}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_193 = core__GEN_183;
  assign _GEN_942 = {_GEN_941,profilePin_193}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_194 = core__GEN_184_0;
  assign _GEN_943 = {_GEN_942,profilePin_194}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_195 = core__GEN_185;
  assign _GEN_944 = {_GEN_943,profilePin_195}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_196 = core__GEN_186;
  assign _GEN_945 = {_GEN_944,profilePin_196}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_197 = core__GEN_187_0;
  assign _GEN_946 = {_GEN_945,profilePin_197}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_198 = core__GEN_188;
  assign _GEN_947 = {_GEN_946,profilePin_198}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_199 = core__GEN_189;
  assign _GEN_948 = {_GEN_947,profilePin_199}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_200 = core__GEN_190;
  assign _GEN_949 = {_GEN_948,profilePin_200}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_201 = core__GEN_191_0;
  assign _GEN_950 = {_GEN_949,profilePin_201}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_202 = core__GEN_192;
  assign _GEN_951 = {_GEN_950,profilePin_202}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_203 = core__GEN_193;
  assign _GEN_952 = {_GEN_951,profilePin_203}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_204 = core__GEN_194_0;
  assign _GEN_953 = {_GEN_952,profilePin_204}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_205 = core__GEN_195;
  assign _GEN_954 = {_GEN_953,profilePin_205}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_206 = core__GEN_196;
  assign _GEN_955 = {_GEN_954,profilePin_206}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_207 = core__GEN_197_0;
  assign _GEN_956 = {_GEN_955,profilePin_207}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_208 = core__GEN_198;
  assign _GEN_957 = {_GEN_956,profilePin_208}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_209 = core__GEN_199;
  assign _GEN_958 = {_GEN_957,profilePin_209}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_210 = core__GEN_200_0;
  assign _GEN_959 = {_GEN_958,profilePin_210}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_211 = core__GEN_201;
  assign _GEN_960 = {_GEN_959,profilePin_211}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_212 = core__GEN_202;
  assign _GEN_961 = {_GEN_960,profilePin_212}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_213 = core__GEN_203_0;
  assign _GEN_962 = {_GEN_961,profilePin_213}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_214 = core__GEN_204;
  assign _GEN_963 = {_GEN_962,profilePin_214}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_215 = core__GEN_205;
  assign _GEN_964 = {_GEN_963,profilePin_215}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_216 = core__GEN_206_0;
  assign _GEN_965 = {_GEN_964,profilePin_216}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_217 = core__GEN_207;
  assign _GEN_966 = {_GEN_965,profilePin_217}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_218 = core__GEN_208;
  assign _GEN_967 = {_GEN_966,profilePin_218}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_219 = core__GEN_209;
  assign _GEN_968 = {_GEN_967,profilePin_219}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_220 = core__GEN_210;
  assign _GEN_969 = {_GEN_968,profilePin_220}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_221 = core__GEN_211;
  assign _GEN_970 = {_GEN_969,profilePin_221}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_222 = core__GEN_212_0;
  assign _GEN_971 = {_GEN_970,profilePin_222}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_223 = core__GEN_213;
  assign _GEN_972 = {_GEN_971,profilePin_223}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_224 = core__GEN_214;
  assign _GEN_973 = {_GEN_972,profilePin_224}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_225 = core__GEN_215;
  assign _GEN_974 = {_GEN_973,profilePin_225}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_226 = core__GEN_216;
  assign _GEN_975 = {_GEN_974,profilePin_226}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_227 = core__GEN_217_0;
  assign _GEN_976 = {_GEN_975,profilePin_227}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_228 = core__GEN_218_0;
  assign _GEN_977 = {_GEN_976,profilePin_228}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_229 = core__GEN_219;
  assign _GEN_978 = {_GEN_977,profilePin_229}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_230 = core__GEN_220;
  assign _GEN_979 = {_GEN_978,profilePin_230}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_231 = core__GEN_221;
  assign _GEN_980 = {_GEN_979,profilePin_231}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_232 = core__GEN_222;
  assign _GEN_981 = {_GEN_980,profilePin_232}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_233 = core__GEN_223_0;
  assign _GEN_982 = {_GEN_981,profilePin_233}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_234 = core__GEN_224_0;
  assign _GEN_983 = {_GEN_982,profilePin_234}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_235 = core__GEN_225;
  assign _GEN_984 = {_GEN_983,profilePin_235}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_236 = core__GEN_226;
  assign _GEN_985 = {_GEN_984,profilePin_236}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_237 = core__GEN_227;
  assign _GEN_986 = {_GEN_985,profilePin_237}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_238 = core__GEN_228;
  assign _GEN_987 = {_GEN_986,profilePin_238}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_239 = core__GEN_229;
  assign _GEN_988 = {_GEN_987,profilePin_239}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_240 = core__GEN_230;
  assign _GEN_989 = {_GEN_988,profilePin_240}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_241 = core__GEN_231;
  assign _GEN_990 = {_GEN_989,profilePin_241}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_242 = core__GEN_232;
  assign _GEN_991 = {_GEN_990,profilePin_242}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_243 = core__GEN_233;
  assign _GEN_992 = {_GEN_991,profilePin_243}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_244 = core__GEN_234;
  assign _GEN_993 = {_GEN_992,profilePin_244}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_245 = core__GEN_235_0;
  assign _GEN_994 = {_GEN_993,profilePin_245}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_246 = core__GEN_236;
  assign _GEN_995 = {_GEN_994,profilePin_246}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_247 = core__GEN_237;
  assign _GEN_996 = {_GEN_995,profilePin_247}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_248 = core__GEN_238_0;
  assign _GEN_997 = {_GEN_996,profilePin_248}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_249 = core__GEN_239_0;
  assign _GEN_998 = {_GEN_997,profilePin_249}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_250 = core__GEN_240;
  assign _GEN_999 = {_GEN_998,profilePin_250}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_251 = core__GEN_241_0;
  assign _GEN_1000 = {_GEN_999,profilePin_251}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_252 = core__GEN_242;
  assign _GEN_1001 = {_GEN_1000,profilePin_252}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_253 = core__GEN_243;
  assign _GEN_1002 = {_GEN_1001,profilePin_253}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_254 = core__GEN_244_0;
  assign _GEN_1003 = {_GEN_1002,profilePin_254}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_255 = core__GEN_245;
  assign _GEN_1004 = {_GEN_1003,profilePin_255}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_256 = core__GEN_246;
  assign _GEN_1005 = {_GEN_1004,profilePin_256}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_257 = core__GEN_247;
  assign _GEN_1006 = {_GEN_1005,profilePin_257}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_258 = core__GEN_248;
  assign _GEN_1007 = {_GEN_1006,profilePin_258}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_259 = core__GEN_249;
  assign _GEN_1008 = {_GEN_1007,profilePin_259}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_260 = core__GEN_250_0;
  assign _GEN_1009 = {_GEN_1008,profilePin_260}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_261 = core__GEN_251;
  assign _GEN_1010 = {_GEN_1009,profilePin_261}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_262 = core__GEN_252;
  assign _GEN_1011 = {_GEN_1010,profilePin_262}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_263 = core__GEN_253_0;
  assign _GEN_1012 = {_GEN_1011,profilePin_263}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_264 = core__GEN_254;
  assign _GEN_1013 = {_GEN_1012,profilePin_264}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_265 = core__GEN_255;
  assign _GEN_1014 = {_GEN_1013,profilePin_265}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_266 = core__GEN_256_0;
  assign _GEN_1015 = {_GEN_1014,profilePin_266}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_267 = core__GEN_257;
  assign _GEN_1016 = {_GEN_1015,profilePin_267}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_268 = core__GEN_258;
  assign _GEN_1017 = {_GEN_1016,profilePin_268}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_269 = core__GEN_259_0;
  assign _GEN_1018 = {_GEN_1017,profilePin_269}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_270 = core__GEN_260;
  assign _GEN_1019 = {_GEN_1018,profilePin_270}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_271 = core__GEN_261;
  assign _GEN_1020 = {_GEN_1019,profilePin_271}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_272 = core__GEN_262_0;
  assign _GEN_1021 = {_GEN_1020,profilePin_272}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_273 = core__GEN_263;
  assign _GEN_1022 = {_GEN_1021,profilePin_273}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_274 = core__GEN_264;
  assign _GEN_1023 = {_GEN_1022,profilePin_274}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_275 = core__GEN_265_0;
  assign _GEN_1024 = {_GEN_1023,profilePin_275}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_276 = core__GEN_266;
  assign _GEN_1025 = {_GEN_1024,profilePin_276}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_277 = core__GEN_267;
  assign _GEN_1026 = {_GEN_1025,profilePin_277}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_278 = core__GEN_268_0;
  assign _GEN_1027 = {_GEN_1026,profilePin_278}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_279 = core__GEN_269;
  assign _GEN_1028 = {_GEN_1027,profilePin_279}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_280 = core__GEN_270;
  assign _GEN_1029 = {_GEN_1028,profilePin_280}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_281 = core__GEN_271_0;
  assign _GEN_1030 = {_GEN_1029,profilePin_281}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_282 = core__GEN_272;
  assign _GEN_1031 = {_GEN_1030,profilePin_282}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_283 = core__GEN_273;
  assign _GEN_1032 = {_GEN_1031,profilePin_283}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_284 = core__GEN_274_0;
  assign _GEN_1033 = {_GEN_1032,profilePin_284}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_285 = core__GEN_275;
  assign _GEN_1034 = {_GEN_1033,profilePin_285}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_286 = core__GEN_276;
  assign _GEN_1035 = {_GEN_1034,profilePin_286}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_287 = core__GEN_277_0;
  assign _GEN_1036 = {_GEN_1035,profilePin_287}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_288 = core__GEN_278;
  assign _GEN_1037 = {_GEN_1036,profilePin_288}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_289 = core__GEN_279;
  assign _GEN_1038 = {_GEN_1037,profilePin_289}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_290 = core__GEN_280_0;
  assign _GEN_1039 = {_GEN_1038,profilePin_290}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_291 = core__GEN_281;
  assign _GEN_1040 = {_GEN_1039,profilePin_291}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_292 = core__GEN_282;
  assign _GEN_1041 = {_GEN_1040,profilePin_292}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_293 = core__GEN_283_0;
  assign _GEN_1042 = {_GEN_1041,profilePin_293}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_294 = core__GEN_284;
  assign _GEN_1043 = {_GEN_1042,profilePin_294}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_295 = core__GEN_285;
  assign _GEN_1044 = {_GEN_1043,profilePin_295}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_296 = core__GEN_286_0;
  assign _GEN_1045 = {_GEN_1044,profilePin_296}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_297 = core__GEN_287;
  assign _GEN_1046 = {_GEN_1045,profilePin_297}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_298 = core__GEN_288;
  assign _GEN_1047 = {_GEN_1046,profilePin_298}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_299 = core__GEN_289_0;
  assign _GEN_1048 = {_GEN_1047,profilePin_299}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_300 = core__GEN_290_0;
  assign _GEN_1049 = {_GEN_1048,profilePin_300}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_301 = core__GEN_291;
  assign _GEN_1050 = {_GEN_1049,profilePin_301}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_302 = core__GEN_292;
  assign _GEN_1051 = {_GEN_1050,profilePin_302}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_303 = core__GEN_293_0;
  assign _GEN_1052 = {_GEN_1051,profilePin_303}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_304 = core__GEN_294;
  assign _GEN_1053 = {_GEN_1052,profilePin_304}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_305 = core__GEN_295;
  assign _GEN_1054 = {_GEN_1053,profilePin_305}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_306 = core__GEN_296_0;
  assign _GEN_1055 = {_GEN_1054,profilePin_306}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_307 = core__GEN_297;
  assign _GEN_1056 = {_GEN_1055,profilePin_307}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_308 = core__GEN_298;
  assign _GEN_1057 = {_GEN_1056,profilePin_308}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_309 = core__GEN_299_0;
  assign _GEN_1058 = {_GEN_1057,profilePin_309}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_310 = core__GEN_300;
  assign _GEN_1059 = {_GEN_1058,profilePin_310}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_311 = core__GEN_301;
  assign _GEN_1060 = {_GEN_1059,profilePin_311}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_312 = core__GEN_302_0;
  assign _GEN_1061 = {_GEN_1060,profilePin_312}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_313 = core__GEN_303;
  assign _GEN_1062 = {_GEN_1061,profilePin_313}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_314 = core__GEN_304;
  assign _GEN_1063 = {_GEN_1062,profilePin_314}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_315 = core__GEN_305_0;
  assign _GEN_1064 = {_GEN_1063,profilePin_315}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_316 = core__GEN_306;
  assign _GEN_1065 = {_GEN_1064,profilePin_316}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_317 = core__GEN_307;
  assign _GEN_1066 = {_GEN_1065,profilePin_317}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_318 = core__GEN_308;
  assign _GEN_1067 = {_GEN_1066,profilePin_318}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_319 = core__GEN_309;
  assign _GEN_1068 = {_GEN_1067,profilePin_319}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_320 = core__GEN_310;
  assign _GEN_1069 = {_GEN_1068,profilePin_320}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_321 = core__GEN_311_0;
  assign _GEN_1070 = {_GEN_1069,profilePin_321}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_322 = core__GEN_312;
  assign _GEN_1071 = {_GEN_1070,profilePin_322}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_323 = core__GEN_313;
  assign _GEN_1072 = {_GEN_1071,profilePin_323}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_324 = core__GEN_314;
  assign _GEN_1073 = {_GEN_1072,profilePin_324}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_325 = core__GEN_315;
  assign _GEN_1074 = {_GEN_1073,profilePin_325}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_326 = core__GEN_316_0;
  assign _GEN_1075 = {_GEN_1074,profilePin_326}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_327 = core__GEN_317_0;
  assign _GEN_1076 = {_GEN_1075,profilePin_327}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_328 = core__GEN_318;
  assign _GEN_1077 = {_GEN_1076,profilePin_328}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_329 = core__GEN_319;
  assign _GEN_1078 = {_GEN_1077,profilePin_329}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_330 = core__GEN_320_0;
  assign _GEN_1079 = {_GEN_1078,profilePin_330}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_331 = core__GEN_321;
  assign _GEN_1080 = {_GEN_1079,profilePin_331}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_332 = core__GEN_322_0;
  assign _GEN_1081 = {_GEN_1080,profilePin_332}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_333 = core__GEN_323_0;
  assign _GEN_1082 = {_GEN_1081,profilePin_333}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_334 = core__GEN_324;
  assign _GEN_1083 = {_GEN_1082,profilePin_334}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_335 = core__GEN_325;
  assign _GEN_1084 = {_GEN_1083,profilePin_335}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_336 = core__GEN_326;
  assign _GEN_1085 = {_GEN_1084,profilePin_336}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_337 = core__GEN_327;
  assign _GEN_1086 = {_GEN_1085,profilePin_337}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_338 = core__GEN_328_0;
  assign _GEN_1087 = {_GEN_1086,profilePin_338}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_339 = core__GEN_329;
  assign _GEN_1088 = {_GEN_1087,profilePin_339}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_340 = core__GEN_330;
  assign _GEN_1089 = {_GEN_1088,profilePin_340}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_341 = core__GEN_331;
  assign _GEN_1090 = {_GEN_1089,profilePin_341}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_342 = core__GEN_332;
  assign _GEN_1091 = {_GEN_1090,profilePin_342}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_343 = core__GEN_333;
  assign _GEN_1092 = {_GEN_1091,profilePin_343}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_344 = core__GEN_334_0;
  assign _GEN_1093 = {_GEN_1092,profilePin_344}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_345 = core__GEN_335;
  assign _GEN_1094 = {_GEN_1093,profilePin_345}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_346 = core__GEN_336;
  assign _GEN_1095 = {_GEN_1094,profilePin_346}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_347 = core__GEN_337_0;
  assign _GEN_1096 = {_GEN_1095,profilePin_347}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_348 = core__GEN_338_0;
  assign _GEN_1097 = {_GEN_1096,profilePin_348}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_349 = core__GEN_339;
  assign _GEN_1098 = {_GEN_1097,profilePin_349}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_350 = core__GEN_340_0;
  assign _GEN_1099 = {_GEN_1098,profilePin_350}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_351 = core__GEN_341;
  assign _GEN_1100 = {_GEN_1099,profilePin_351}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_352 = core__GEN_342;
  assign _GEN_1101 = {_GEN_1100,profilePin_352}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_353 = core__GEN_343_0;
  assign _GEN_1102 = {_GEN_1101,profilePin_353}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_354 = core__GEN_344;
  assign _GEN_1103 = {_GEN_1102,profilePin_354}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_355 = core__GEN_345;
  assign _GEN_1104 = {_GEN_1103,profilePin_355}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_356 = core__GEN_346_0;
  assign _GEN_1105 = {_GEN_1104,profilePin_356}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_357 = core__GEN_347;
  assign _GEN_1106 = {_GEN_1105,profilePin_357}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_358 = core__GEN_348;
  assign _GEN_1107 = {_GEN_1106,profilePin_358}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_359 = core__GEN_349_0;
  assign _GEN_1108 = {_GEN_1107,profilePin_359}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_360 = core__GEN_350;
  assign _GEN_1109 = {_GEN_1108,profilePin_360}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_361 = core__GEN_351;
  assign _GEN_1110 = {_GEN_1109,profilePin_361}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_362 = core__GEN_352_0;
  assign _GEN_1111 = {_GEN_1110,profilePin_362}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_363 = core__GEN_353;
  assign _GEN_1112 = {_GEN_1111,profilePin_363}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_364 = core__GEN_354;
  assign _GEN_1113 = {_GEN_1112,profilePin_364}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_365 = core__GEN_355_0;
  assign _GEN_1114 = {_GEN_1113,profilePin_365}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_366 = core__GEN_356;
  assign _GEN_1115 = {_GEN_1114,profilePin_366}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_367 = core__GEN_357;
  assign _GEN_1116 = {_GEN_1115,profilePin_367}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_368 = core__GEN_358_0;
  assign _GEN_1117 = {_GEN_1116,profilePin_368}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_369 = core__GEN_359;
  assign _GEN_1118 = {_GEN_1117,profilePin_369}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_370 = core__GEN_360;
  assign _GEN_1119 = {_GEN_1118,profilePin_370}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_371 = core__GEN_361_0;
  assign _GEN_1120 = {_GEN_1119,profilePin_371}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_372 = core__GEN_362;
  assign _GEN_1121 = {_GEN_1120,profilePin_372}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_373 = core__GEN_363;
  assign _GEN_1122 = {_GEN_1121,profilePin_373}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_374 = core__GEN_364_0;
  assign _GEN_1123 = {_GEN_1122,profilePin_374}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_375 = core__GEN_365;
  assign _GEN_1124 = {_GEN_1123,profilePin_375}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_376 = core__GEN_366;
  assign _GEN_1125 = {_GEN_1124,profilePin_376}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_377 = core__GEN_367_0;
  assign _GEN_1126 = {_GEN_1125,profilePin_377}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_378 = core__GEN_368;
  assign _GEN_1127 = {_GEN_1126,profilePin_378}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_379 = core__GEN_369;
  assign _GEN_1128 = {_GEN_1127,profilePin_379}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_380 = core__GEN_370_0;
  assign _GEN_1129 = {_GEN_1128,profilePin_380}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_381 = core__GEN_371;
  assign _GEN_1130 = {_GEN_1129,profilePin_381}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_382 = core__GEN_372;
  assign _GEN_1131 = {_GEN_1130,profilePin_382}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_383 = core__GEN_373_0;
  assign _GEN_1132 = {_GEN_1131,profilePin_383}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_384 = core__GEN_374;
  assign _GEN_1133 = {_GEN_1132,profilePin_384}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_385 = core__GEN_375;
  assign _GEN_1134 = {_GEN_1133,profilePin_385}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_386 = core__GEN_376_0;
  assign _GEN_1135 = {_GEN_1134,profilePin_386}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_387 = core__GEN_377;
  assign _GEN_1136 = {_GEN_1135,profilePin_387}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_388 = core__GEN_378;
  assign _GEN_1137 = {_GEN_1136,profilePin_388}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_389 = core__GEN_379_0;
  assign _GEN_1138 = {_GEN_1137,profilePin_389}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_390 = core__GEN_380;
  assign _GEN_1139 = {_GEN_1138,profilePin_390}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_391 = core__GEN_381;
  assign _GEN_1140 = {_GEN_1139,profilePin_391}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_392 = core__GEN_382_0;
  assign _GEN_1141 = {_GEN_1140,profilePin_392}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_393 = core__GEN_383;
  assign _GEN_1142 = {_GEN_1141,profilePin_393}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_394 = core__GEN_384;
  assign _GEN_1143 = {_GEN_1142,profilePin_394}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_395 = core__GEN_385_0;
  assign _GEN_1144 = {_GEN_1143,profilePin_395}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_396 = core__GEN_386;
  assign _GEN_1145 = {_GEN_1144,profilePin_396}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_397 = core__GEN_387;
  assign _GEN_1146 = {_GEN_1145,profilePin_397}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_398 = core__GEN_388_0;
  assign _GEN_1147 = {_GEN_1146,profilePin_398}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_399 = core__GEN_389;
  assign _GEN_1148 = {_GEN_1147,profilePin_399}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_400 = core__GEN_390;
  assign _GEN_1149 = {_GEN_1148,profilePin_400}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_401 = core__GEN_391;
  assign _GEN_1150 = {_GEN_1149,profilePin_401}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_402 = core__GEN_392;
  assign _GEN_1151 = {_GEN_1150,profilePin_402}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_403 = core__GEN_393;
  assign _GEN_1152 = {_GEN_1151,profilePin_403}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_404 = core__GEN_394;
  assign _GEN_1153 = {_GEN_1152,profilePin_404}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_405 = core__GEN_395;
  assign _GEN_1154 = {_GEN_1153,profilePin_405}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_406 = core__GEN_396;
  assign _GEN_1155 = {_GEN_1154,profilePin_406}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_407 = core__GEN_397;
  assign _GEN_1156 = {_GEN_1155,profilePin_407}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_408 = core__GEN_398;
  assign _GEN_1157 = {_GEN_1156,profilePin_408}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_409 = core__GEN_399;
  assign _GEN_1158 = {_GEN_1157,profilePin_409}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_410 = core__GEN_400;
  assign _GEN_1159 = {_GEN_1158,profilePin_410}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_411 = core__GEN_401;
  assign _GEN_1160 = {_GEN_1159,profilePin_411}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_412 = core__GEN_402;
  assign _GEN_1161 = {_GEN_1160,profilePin_412}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_413 = core__GEN_403;
  assign _GEN_1162 = {_GEN_1161,profilePin_413}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_414 = core__GEN_404;
  assign _GEN_1163 = {_GEN_1162,profilePin_414}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_415 = core__GEN_405;
  assign _GEN_1164 = {_GEN_1163,profilePin_415}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_416 = core__GEN_406;
  assign _GEN_1165 = {_GEN_1164,profilePin_416}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_417 = core__GEN_407;
  assign _GEN_1166 = {_GEN_1165,profilePin_417}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_418 = core__GEN_408;
  assign _GEN_1167 = {_GEN_1166,profilePin_418}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_419 = core__GEN_409;
  assign _GEN_1168 = {_GEN_1167,profilePin_419}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_420 = core__GEN_410;
  assign _GEN_1169 = {_GEN_1168,profilePin_420}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_421 = core__GEN_411;
  assign _GEN_1170 = {_GEN_1169,profilePin_421}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_422 = core__GEN_412;
  assign _GEN_1171 = {_GEN_1170,profilePin_422}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_423 = core__GEN_413;
  assign _GEN_1172 = {_GEN_1171,profilePin_423}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_424 = core__GEN_414;
  assign _GEN_1173 = {_GEN_1172,profilePin_424}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_425 = core__GEN_415;
  assign _GEN_1174 = {_GEN_1173,profilePin_425}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_426 = core__GEN_416;
  assign _GEN_1175 = {_GEN_1174,profilePin_426}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_427 = core__GEN_417;
  assign _GEN_1176 = {_GEN_1175,profilePin_427}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_428 = core__GEN_418;
  assign _GEN_1177 = {_GEN_1176,profilePin_428}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_429 = core__GEN_419;
  assign _GEN_1178 = {_GEN_1177,profilePin_429}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_430 = core__GEN_420;
  assign _GEN_1179 = {_GEN_1178,profilePin_430}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_431 = core__GEN_421;
  assign _GEN_1180 = {_GEN_1179,profilePin_431}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_432 = core__GEN_422;
  assign _GEN_1181 = {_GEN_1180,profilePin_432}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_433 = core__GEN_423;
  assign _GEN_1182 = {_GEN_1181,profilePin_433}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_434 = core__GEN_424;
  assign _GEN_1183 = {_GEN_1182,profilePin_434}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_435 = core__GEN_425;
  assign _GEN_1184 = {_GEN_1183,profilePin_435}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_436 = core__GEN_426;
  assign _GEN_1185 = {_GEN_1184,profilePin_436}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_437 = core__GEN_427;
  assign _GEN_1186 = {_GEN_1185,profilePin_437}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_438 = core__GEN_428;
  assign _GEN_1187 = {_GEN_1186,profilePin_438}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_439 = core__GEN_429;
  assign _GEN_1188 = {_GEN_1187,profilePin_439}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_440 = core__GEN_0;
  assign _GEN_1189 = {_GEN_1188,profilePin_440}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_441 = core__GEN_1_3;
  assign _GEN_1190 = {_GEN_1189,profilePin_441}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_442 = core__GEN_2;
  assign _GEN_1191 = {_GEN_1190,profilePin_442}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_443 = core__GEN_3_4;
  assign _GEN_1192 = {_GEN_1191,profilePin_443}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_444 = core__GEN_4_1;
  assign _GEN_1193 = {_GEN_1192,profilePin_444}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_445 = core__GEN_5_0;
  assign _GEN_1194 = {_GEN_1193,profilePin_445}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_446 = core__GEN_6_4;
  assign _GEN_1195 = {_GEN_1194,profilePin_446}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_447 = core__GEN_7_1;
  assign _GEN_1196 = {_GEN_1195,profilePin_447}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_448 = core__GEN_8;
  assign _GEN_1197 = {_GEN_1196,profilePin_448}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_449 = core__GEN_9_0;
  assign _GEN_1198 = {_GEN_1197,profilePin_449}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_450 = core__GEN_10_0;
  assign _GEN_1199 = {_GEN_1198,profilePin_450}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_451 = core__GEN_3_2;
  assign _GEN_1200 = {_GEN_1199,profilePin_451}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_452 = core__GEN_5_4;
  assign _GEN_1201 = {_GEN_1200,profilePin_452}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_453 = core__GEN_7_2;
  assign _GEN_1202 = {_GEN_1201,profilePin_453}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_454 = core__GEN_11;
  assign _GEN_1203 = {_GEN_1202,profilePin_454}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_455 = core__GEN_15_1;
  assign _GEN_1204 = {_GEN_1203,profilePin_455}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_456 = core__GEN_146_0;
  assign _GEN_1205 = {_GEN_1204,profilePin_456}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_457 = core__GEN_147_0;
  assign _GEN_1206 = {_GEN_1205,profilePin_457}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_458 = core__GEN_149_0;
  assign _GEN_1207 = {_GEN_1206,profilePin_458}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_459 = core__GEN_150_0;
  assign _GEN_1208 = {_GEN_1207,profilePin_459}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_460 = core__GEN_151;
  assign _GEN_1209 = {_GEN_1208,profilePin_460}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_461 = core__GEN_152_0;
  assign _GEN_1210 = {_GEN_1209,profilePin_461}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_462 = core__GEN_153_0;
  assign _GEN_1211 = {_GEN_1210,profilePin_462}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_463 = core__GEN_154;
  assign _GEN_1212 = {_GEN_1211,profilePin_463}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_464 = core__GEN_155_0;
  assign _GEN_1213 = {_GEN_1212,profilePin_464}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_465 = core__GEN_156_0;
  assign _GEN_1214 = {_GEN_1213,profilePin_465}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_466 = core__GEN_157;
  assign _GEN_1215 = {_GEN_1214,profilePin_466}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_467 = core__GEN_158_0;
  assign _GEN_1216 = {_GEN_1215,profilePin_467}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_468 = core__GEN_159_0;
  assign _GEN_1217 = {_GEN_1216,profilePin_468}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_469 = core__GEN_160;
  assign _GEN_1218 = {_GEN_1217,profilePin_469}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_470 = core__GEN_161_0;
  assign _GEN_1219 = {_GEN_1218,profilePin_470}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_471 = core__GEN_162_0;
  assign _GEN_1220 = {_GEN_1219,profilePin_471}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_472 = core__GEN_163;
  assign _GEN_1221 = {_GEN_1220,profilePin_472}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_473 = core__GEN_164_0;
  assign _GEN_1222 = {_GEN_1221,profilePin_473}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_474 = core__GEN_165_0;
  assign _GEN_1223 = {_GEN_1222,profilePin_474}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_475 = core__GEN_166;
  assign _GEN_1224 = {_GEN_1223,profilePin_475}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_476 = core__GEN_167_0;
  assign _GEN_1225 = {_GEN_1224,profilePin_476}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_477 = core__GEN_168_0;
  assign _GEN_1226 = {_GEN_1225,profilePin_477}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_478 = core__GEN_169;
  assign _GEN_1227 = {_GEN_1226,profilePin_478}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_479 = core__GEN_170_0;
  assign _GEN_1228 = {_GEN_1227,profilePin_479}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_480 = core__GEN_171_0;
  assign _GEN_1229 = {_GEN_1228,profilePin_480}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_481 = core__GEN_172;
  assign _GEN_1230 = {_GEN_1229,profilePin_481}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_482 = core__GEN_173_0;
  assign _GEN_1231 = {_GEN_1230,profilePin_482}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_483 = core__GEN_174_0;
  assign _GEN_1232 = {_GEN_1231,profilePin_483}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_484 = core__GEN_175;
  assign _GEN_1233 = {_GEN_1232,profilePin_484}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_485 = core__GEN_176_0;
  assign _GEN_1234 = {_GEN_1233,profilePin_485}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_486 = core__GEN_177_0;
  assign _GEN_1235 = {_GEN_1234,profilePin_486}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_487 = core__GEN_178;
  assign _GEN_1236 = {_GEN_1235,profilePin_487}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_488 = core__GEN_179_0;
  assign _GEN_1237 = {_GEN_1236,profilePin_488}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_489 = core__GEN_180_0;
  assign _GEN_1238 = {_GEN_1237,profilePin_489}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_490 = core__GEN_181;
  assign _GEN_1239 = {_GEN_1238,profilePin_490}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_491 = core__GEN_182_0;
  assign _GEN_1240 = {_GEN_1239,profilePin_491}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_492 = core__GEN_183_0;
  assign _GEN_1241 = {_GEN_1240,profilePin_492}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_493 = core__GEN_184;
  assign _GEN_1242 = {_GEN_1241,profilePin_493}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_494 = core__GEN_185_0;
  assign _GEN_1243 = {_GEN_1242,profilePin_494}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_495 = core__GEN_186_0;
  assign _GEN_1244 = {_GEN_1243,profilePin_495}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_496 = core__GEN_187;
  assign _GEN_1245 = {_GEN_1244,profilePin_496}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_497 = core__GEN_188_0;
  assign _GEN_1246 = {_GEN_1245,profilePin_497}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_498 = core__GEN_189_0;
  assign _GEN_1247 = {_GEN_1246,profilePin_498}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_499 = core__GEN_190_0;
  assign _GEN_1248 = {_GEN_1247,profilePin_499}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_500 = core__GEN_191;
  assign _GEN_1249 = {_GEN_1248,profilePin_500}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_501 = core__GEN_192_0;
  assign _GEN_1250 = {_GEN_1249,profilePin_501}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_502 = core__GEN_193_0;
  assign _GEN_1251 = {_GEN_1250,profilePin_502}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_503 = core__GEN_194;
  assign _GEN_1252 = {_GEN_1251,profilePin_503}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_504 = core__GEN_195_0;
  assign _GEN_1253 = {_GEN_1252,profilePin_504}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_505 = core__GEN_196_0;
  assign _GEN_1254 = {_GEN_1253,profilePin_505}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_506 = core__GEN_197;
  assign _GEN_1255 = {_GEN_1254,profilePin_506}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_507 = core__GEN_198_0;
  assign _GEN_1256 = {_GEN_1255,profilePin_507}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_508 = core__GEN_199_0;
  assign _GEN_1257 = {_GEN_1256,profilePin_508}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_509 = core__GEN_200;
  assign _GEN_1258 = {_GEN_1257,profilePin_509}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_510 = core__GEN_201_0;
  assign _GEN_1259 = {_GEN_1258,profilePin_510}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_511 = core__GEN_202_0;
  assign _GEN_1260 = {_GEN_1259,profilePin_511}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_512 = core__GEN_203;
  assign _GEN_1261 = {_GEN_1260,profilePin_512}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_513 = core__GEN_204_0;
  assign _GEN_1262 = {_GEN_1261,profilePin_513}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_514 = core__GEN_205_0;
  assign _GEN_1263 = {_GEN_1262,profilePin_514}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_515 = core__GEN_206;
  assign _GEN_1264 = {_GEN_1263,profilePin_515}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_516 = core__GEN_207_0;
  assign _GEN_1265 = {_GEN_1264,profilePin_516}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_517 = core__GEN_208_0;
  assign _GEN_1266 = {_GEN_1265,profilePin_517}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_518 = core__GEN_209_0;
  assign _GEN_1267 = {_GEN_1266,profilePin_518}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_519 = core__GEN_210_0;
  assign _GEN_1268 = {_GEN_1267,profilePin_519}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_520 = core__GEN_211_0;
  assign _GEN_1269 = {_GEN_1268,profilePin_520}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_521 = core__GEN_212;
  assign _GEN_1270 = {_GEN_1269,profilePin_521}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_522 = core__GEN_213_0;
  assign _GEN_1271 = {_GEN_1270,profilePin_522}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_523 = core__GEN_214_0;
  assign _GEN_1272 = {_GEN_1271,profilePin_523}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_524 = core__GEN_215_0;
  assign _GEN_1273 = {_GEN_1272,profilePin_524}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_525 = core__GEN_216_0;
  assign _GEN_1274 = {_GEN_1273,profilePin_525}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_526 = core__GEN_217;
  assign _GEN_1275 = {_GEN_1274,profilePin_526}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_527 = core__GEN_218;
  assign _GEN_1276 = {_GEN_1275,profilePin_527}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_528 = core__GEN_219_0;
  assign _GEN_1277 = {_GEN_1276,profilePin_528}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_529 = core__GEN_220_0;
  assign _GEN_1278 = {_GEN_1277,profilePin_529}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_530 = core__GEN_221_0;
  assign _GEN_1279 = {_GEN_1278,profilePin_530}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_531 = core__GEN_222_0;
  assign _GEN_1280 = {_GEN_1279,profilePin_531}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_532 = core__GEN_223;
  assign _GEN_1281 = {_GEN_1280,profilePin_532}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_533 = core__GEN_224;
  assign _GEN_1282 = {_GEN_1281,profilePin_533}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_534 = core__GEN_225_0;
  assign _GEN_1283 = {_GEN_1282,profilePin_534}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_535 = core__GEN_226_0;
  assign _GEN_1284 = {_GEN_1283,profilePin_535}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_536 = core__GEN_227_0;
  assign _GEN_1285 = {_GEN_1284,profilePin_536}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_537 = core__GEN_228_0;
  assign _GEN_1286 = {_GEN_1285,profilePin_537}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_538 = core__GEN_229_0;
  assign _GEN_1287 = {_GEN_1286,profilePin_538}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_539 = core__GEN_230_0;
  assign _GEN_1288 = {_GEN_1287,profilePin_539}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_540 = core__GEN_231_0;
  assign _GEN_1289 = {_GEN_1288,profilePin_540}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_541 = core__GEN_232_0;
  assign _GEN_1290 = {_GEN_1289,profilePin_541}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_542 = core__GEN_233_0;
  assign _GEN_1291 = {_GEN_1290,profilePin_542}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_543 = core__GEN_234_0;
  assign _GEN_1292 = {_GEN_1291,profilePin_543}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_544 = core__GEN_235;
  assign _GEN_1293 = {_GEN_1292,profilePin_544}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_545 = core__GEN_236_0;
  assign _GEN_1294 = {_GEN_1293,profilePin_545}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_546 = core__GEN_237_0;
  assign _GEN_1295 = {_GEN_1294,profilePin_546}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_547 = core__GEN_238;
  assign _GEN_1296 = {_GEN_1295,profilePin_547}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_548 = core__GEN_239;
  assign _GEN_1297 = {_GEN_1296,profilePin_548}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_549 = core__GEN_240_0;
  assign _GEN_1298 = {_GEN_1297,profilePin_549}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_550 = core__GEN_241;
  assign _GEN_1299 = {_GEN_1298,profilePin_550}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_551 = core__GEN_242_0;
  assign _GEN_1300 = {_GEN_1299,profilePin_551}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_552 = core__GEN_243_0;
  assign _GEN_1301 = {_GEN_1300,profilePin_552}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_553 = core__GEN_244;
  assign _GEN_1302 = {_GEN_1301,profilePin_553}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_554 = core__GEN_245_0;
  assign _GEN_1303 = {_GEN_1302,profilePin_554}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_555 = core__GEN_246_0;
  assign _GEN_1304 = {_GEN_1303,profilePin_555}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_556 = core__GEN_247_0;
  assign _GEN_1305 = {_GEN_1304,profilePin_556}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_557 = core__GEN_248_0;
  assign _GEN_1306 = {_GEN_1305,profilePin_557}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_558 = core__GEN_249_0;
  assign _GEN_1307 = {_GEN_1306,profilePin_558}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_559 = core__GEN_250;
  assign _GEN_1308 = {_GEN_1307,profilePin_559}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_560 = core__GEN_251_0;
  assign _GEN_1309 = {_GEN_1308,profilePin_560}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_561 = core__GEN_252_0;
  assign _GEN_1310 = {_GEN_1309,profilePin_561}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_562 = core__GEN_253;
  assign _GEN_1311 = {_GEN_1310,profilePin_562}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_563 = core__GEN_254_0;
  assign _GEN_1312 = {_GEN_1311,profilePin_563}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_564 = core__GEN_255_0;
  assign _GEN_1313 = {_GEN_1312,profilePin_564}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_565 = core__GEN_256;
  assign _GEN_1314 = {_GEN_1313,profilePin_565}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_566 = core__GEN_257_0;
  assign _GEN_1315 = {_GEN_1314,profilePin_566}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_567 = core__GEN_258_0;
  assign _GEN_1316 = {_GEN_1315,profilePin_567}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_568 = core__GEN_259;
  assign _GEN_1317 = {_GEN_1316,profilePin_568}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_569 = core__GEN_260_0;
  assign _GEN_1318 = {_GEN_1317,profilePin_569}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_570 = core__GEN_261_0;
  assign _GEN_1319 = {_GEN_1318,profilePin_570}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_571 = core__GEN_262;
  assign _GEN_1320 = {_GEN_1319,profilePin_571}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_572 = core__GEN_263_0;
  assign _GEN_1321 = {_GEN_1320,profilePin_572}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_573 = core__GEN_264_0;
  assign _GEN_1322 = {_GEN_1321,profilePin_573}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_574 = core__GEN_265;
  assign _GEN_1323 = {_GEN_1322,profilePin_574}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_575 = core__GEN_266_0;
  assign _GEN_1324 = {_GEN_1323,profilePin_575}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_576 = core__GEN_267_0;
  assign _GEN_1325 = {_GEN_1324,profilePin_576}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_577 = core__GEN_268;
  assign _GEN_1326 = {_GEN_1325,profilePin_577}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_578 = core__GEN_269_0;
  assign _GEN_1327 = {_GEN_1326,profilePin_578}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_579 = core__GEN_270_0;
  assign _GEN_1328 = {_GEN_1327,profilePin_579}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_580 = core__GEN_271;
  assign _GEN_1329 = {_GEN_1328,profilePin_580}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_581 = core__GEN_272_0;
  assign _GEN_1330 = {_GEN_1329,profilePin_581}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_582 = core__GEN_273_0;
  assign _GEN_1331 = {_GEN_1330,profilePin_582}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_583 = core__GEN_274;
  assign _GEN_1332 = {_GEN_1331,profilePin_583}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_584 = core__GEN_275_0;
  assign _GEN_1333 = {_GEN_1332,profilePin_584}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_585 = core__GEN_276_0;
  assign _GEN_1334 = {_GEN_1333,profilePin_585}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_586 = core__GEN_277;
  assign _GEN_1335 = {_GEN_1334,profilePin_586}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_587 = core__GEN_278_0;
  assign _GEN_1336 = {_GEN_1335,profilePin_587}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_588 = core__GEN_279_0;
  assign _GEN_1337 = {_GEN_1336,profilePin_588}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_589 = core__GEN_280;
  assign _GEN_1338 = {_GEN_1337,profilePin_589}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_590 = core__GEN_281_0;
  assign _GEN_1339 = {_GEN_1338,profilePin_590}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_591 = core__GEN_282_0;
  assign _GEN_1340 = {_GEN_1339,profilePin_591}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_592 = core__GEN_283;
  assign _GEN_1341 = {_GEN_1340,profilePin_592}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_593 = core__GEN_284_0;
  assign _GEN_1342 = {_GEN_1341,profilePin_593}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_594 = core__GEN_285_0;
  assign _GEN_1343 = {_GEN_1342,profilePin_594}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_595 = core__GEN_286;
  assign _GEN_1344 = {_GEN_1343,profilePin_595}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_596 = core__GEN_287_0;
  assign _GEN_1345 = {_GEN_1344,profilePin_596}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_597 = core__GEN_288_0;
  assign _GEN_1346 = {_GEN_1345,profilePin_597}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_598 = core__GEN_289;
  assign _GEN_1347 = {_GEN_1346,profilePin_598}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_599 = core__GEN_290;
  assign _GEN_1348 = {_GEN_1347,profilePin_599}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_600 = core__GEN_291_0;
  assign _GEN_1349 = {_GEN_1348,profilePin_600}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_601 = core__GEN_292_0;
  assign _GEN_1350 = {_GEN_1349,profilePin_601}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_602 = core__GEN_293;
  assign _GEN_1351 = {_GEN_1350,profilePin_602}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_603 = core__GEN_294_0;
  assign _GEN_1352 = {_GEN_1351,profilePin_603}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_604 = core__GEN_295_0;
  assign _GEN_1353 = {_GEN_1352,profilePin_604}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_605 = core__GEN_296;
  assign _GEN_1354 = {_GEN_1353,profilePin_605}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_606 = core__GEN_297_0;
  assign _GEN_1355 = {_GEN_1354,profilePin_606}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_607 = core__GEN_298_0;
  assign _GEN_1356 = {_GEN_1355,profilePin_607}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_608 = core__GEN_299;
  assign _GEN_1357 = {_GEN_1356,profilePin_608}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_609 = core__GEN_300_0;
  assign _GEN_1358 = {_GEN_1357,profilePin_609}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_610 = core__GEN_301_0;
  assign _GEN_1359 = {_GEN_1358,profilePin_610}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_611 = core__GEN_302;
  assign _GEN_1360 = {_GEN_1359,profilePin_611}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_612 = core__GEN_303_0;
  assign _GEN_1361 = {_GEN_1360,profilePin_612}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_613 = core__GEN_304_0;
  assign _GEN_1362 = {_GEN_1361,profilePin_613}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_614 = core__GEN_305;
  assign _GEN_1363 = {_GEN_1362,profilePin_614}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_615 = core__GEN_306_0;
  assign _GEN_1364 = {_GEN_1363,profilePin_615}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_616 = core__GEN_307_0;
  assign _GEN_1365 = {_GEN_1364,profilePin_616}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_617 = core__GEN_308_0;
  assign _GEN_1366 = {_GEN_1365,profilePin_617}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_618 = core__GEN_309_0;
  assign _GEN_1367 = {_GEN_1366,profilePin_618}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_619 = core__GEN_310_0;
  assign _GEN_1368 = {_GEN_1367,profilePin_619}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_620 = core__GEN_311;
  assign _GEN_1369 = {_GEN_1368,profilePin_620}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_621 = core__GEN_312_0;
  assign _GEN_1370 = {_GEN_1369,profilePin_621}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_622 = core__GEN_313_0;
  assign _GEN_1371 = {_GEN_1370,profilePin_622}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_623 = core__GEN_314_0;
  assign _GEN_1372 = {_GEN_1371,profilePin_623}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_624 = core__GEN_315_0;
  assign _GEN_1373 = {_GEN_1372,profilePin_624}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_625 = core__GEN_316;
  assign _GEN_1374 = {_GEN_1373,profilePin_625}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_626 = core__GEN_317;
  assign _GEN_1375 = {_GEN_1374,profilePin_626}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_627 = core__GEN_318_0;
  assign _GEN_1376 = {_GEN_1375,profilePin_627}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_628 = core__GEN_319_0;
  assign _GEN_1377 = {_GEN_1376,profilePin_628}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_629 = core__GEN_320;
  assign _GEN_1378 = {_GEN_1377,profilePin_629}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_630 = core__GEN_321_0;
  assign _GEN_1379 = {_GEN_1378,profilePin_630}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_631 = core__GEN_322;
  assign _GEN_1380 = {_GEN_1379,profilePin_631}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_632 = core__GEN_323;
  assign _GEN_1381 = {_GEN_1380,profilePin_632}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_633 = core__GEN_324_0;
  assign _GEN_1382 = {_GEN_1381,profilePin_633}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_634 = core__GEN_325_0;
  assign _GEN_1383 = {_GEN_1382,profilePin_634}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_635 = core__GEN_326_0;
  assign _GEN_1384 = {_GEN_1383,profilePin_635}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_636 = core__GEN_327_0;
  assign _GEN_1385 = {_GEN_1384,profilePin_636}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_637 = core__GEN_328;
  assign _GEN_1386 = {_GEN_1385,profilePin_637}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_638 = core__GEN_329_0;
  assign _GEN_1387 = {_GEN_1386,profilePin_638}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_639 = core__GEN_330_0;
  assign _GEN_1388 = {_GEN_1387,profilePin_639}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_640 = core__GEN_331_0;
  assign _GEN_1389 = {_GEN_1388,profilePin_640}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_641 = core__GEN_332_0;
  assign _GEN_1390 = {_GEN_1389,profilePin_641}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_642 = core__GEN_333_0;
  assign _GEN_1391 = {_GEN_1390,profilePin_642}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_643 = core__GEN_334;
  assign _GEN_1392 = {_GEN_1391,profilePin_643}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_644 = core__GEN_335_0;
  assign _GEN_1393 = {_GEN_1392,profilePin_644}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_645 = core__GEN_336_0;
  assign _GEN_1394 = {_GEN_1393,profilePin_645}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_646 = core__GEN_337;
  assign _GEN_1395 = {_GEN_1394,profilePin_646}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_647 = core__GEN_338;
  assign _GEN_1396 = {_GEN_1395,profilePin_647}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_648 = core__GEN_339_0;
  assign _GEN_1397 = {_GEN_1396,profilePin_648}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_649 = core__GEN_340;
  assign _GEN_1398 = {_GEN_1397,profilePin_649}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_650 = core__GEN_341_0;
  assign _GEN_1399 = {_GEN_1398,profilePin_650}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_651 = core__GEN_342_0;
  assign _GEN_1400 = {_GEN_1399,profilePin_651}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_652 = core__GEN_343;
  assign _GEN_1401 = {_GEN_1400,profilePin_652}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_653 = core__GEN_344_0;
  assign _GEN_1402 = {_GEN_1401,profilePin_653}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_654 = core__GEN_345_0;
  assign _GEN_1403 = {_GEN_1402,profilePin_654}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_655 = core__GEN_346;
  assign _GEN_1404 = {_GEN_1403,profilePin_655}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_656 = core__GEN_347_0;
  assign _GEN_1405 = {_GEN_1404,profilePin_656}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_657 = core__GEN_348_0;
  assign _GEN_1406 = {_GEN_1405,profilePin_657}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_658 = core__GEN_349;
  assign _GEN_1407 = {_GEN_1406,profilePin_658}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_659 = core__GEN_350_0;
  assign _GEN_1408 = {_GEN_1407,profilePin_659}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_660 = core__GEN_351_0;
  assign _GEN_1409 = {_GEN_1408,profilePin_660}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_661 = core__GEN_352;
  assign _GEN_1410 = {_GEN_1409,profilePin_661}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_662 = core__GEN_353_0;
  assign _GEN_1411 = {_GEN_1410,profilePin_662}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_663 = core__GEN_354_0;
  assign _GEN_1412 = {_GEN_1411,profilePin_663}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_664 = core__GEN_355;
  assign _GEN_1413 = {_GEN_1412,profilePin_664}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_665 = core__GEN_356_0;
  assign _GEN_1414 = {_GEN_1413,profilePin_665}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_666 = core__GEN_357_0;
  assign _GEN_1415 = {_GEN_1414,profilePin_666}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_667 = core__GEN_358;
  assign _GEN_1416 = {_GEN_1415,profilePin_667}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_668 = core__GEN_359_0;
  assign _GEN_1417 = {_GEN_1416,profilePin_668}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_669 = core__GEN_360_0;
  assign _GEN_1418 = {_GEN_1417,profilePin_669}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_670 = core__GEN_361;
  assign _GEN_1419 = {_GEN_1418,profilePin_670}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_671 = core__GEN_362_0;
  assign _GEN_1420 = {_GEN_1419,profilePin_671}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_672 = core__GEN_363_0;
  assign _GEN_1421 = {_GEN_1420,profilePin_672}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_673 = core__GEN_364;
  assign _GEN_1422 = {_GEN_1421,profilePin_673}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_674 = core__GEN_365_0;
  assign _GEN_1423 = {_GEN_1422,profilePin_674}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_675 = core__GEN_366_0;
  assign _GEN_1424 = {_GEN_1423,profilePin_675}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_676 = core__GEN_367;
  assign _GEN_1425 = {_GEN_1424,profilePin_676}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_677 = core__GEN_368_0;
  assign _GEN_1426 = {_GEN_1425,profilePin_677}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_678 = core__GEN_369_0;
  assign _GEN_1427 = {_GEN_1426,profilePin_678}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_679 = core__GEN_370;
  assign _GEN_1428 = {_GEN_1427,profilePin_679}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_680 = core__GEN_371_0;
  assign _GEN_1429 = {_GEN_1428,profilePin_680}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_681 = core__GEN_372_0;
  assign _GEN_1430 = {_GEN_1429,profilePin_681}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_682 = core__GEN_373;
  assign _GEN_1431 = {_GEN_1430,profilePin_682}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_683 = core__GEN_374_0;
  assign _GEN_1432 = {_GEN_1431,profilePin_683}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_684 = core__GEN_375_0;
  assign _GEN_1433 = {_GEN_1432,profilePin_684}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_685 = core__GEN_376;
  assign _GEN_1434 = {_GEN_1433,profilePin_685}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_686 = core__GEN_377_0;
  assign _GEN_1435 = {_GEN_1434,profilePin_686}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_687 = core__GEN_378_0;
  assign _GEN_1436 = {_GEN_1435,profilePin_687}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_688 = core__GEN_379;
  assign _GEN_1437 = {_GEN_1436,profilePin_688}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_689 = core__GEN_380_0;
  assign _GEN_1438 = {_GEN_1437,profilePin_689}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_690 = core__GEN_381_0;
  assign _GEN_1439 = {_GEN_1438,profilePin_690}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_691 = core__GEN_382;
  assign _GEN_1440 = {_GEN_1439,profilePin_691}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_692 = core__GEN_383_0;
  assign _GEN_1441 = {_GEN_1440,profilePin_692}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_693 = core__GEN_384_0;
  assign _GEN_1442 = {_GEN_1441,profilePin_693}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_694 = core__GEN_385;
  assign _GEN_1443 = {_GEN_1442,profilePin_694}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_695 = core__GEN_386_0;
  assign _GEN_1444 = {_GEN_1443,profilePin_695}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_696 = core__GEN_387_0;
  assign _GEN_1445 = {_GEN_1444,profilePin_696}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_698 = core__GEN_0_2;
  assign _GEN_1446 = {_GEN_1445,profilePin_698}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_699 = core__GEN_1_1;
  assign _GEN_1447 = {_GEN_1446,profilePin_699}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_700 = core__GEN_2_0;
  assign _GEN_1448 = {_GEN_1447,profilePin_700}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_701 = core__GEN_3_0;
  assign _GEN_1449 = {_GEN_1448,profilePin_701}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_702 = core__GEN_4_2;
  assign _GEN_1450 = {_GEN_1449,profilePin_702}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_703 = core__GEN_5_1;
  assign _GEN_1451 = {_GEN_1450,profilePin_703}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_704 = core__GEN_6;
  assign _GEN_1452 = {_GEN_1451,profilePin_704}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_705 = core__GEN_7_3;
  assign _GEN_1453 = {_GEN_1452,profilePin_705}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_706 = core__GEN_8_1;
  assign _GEN_1454 = {_GEN_1453,profilePin_706}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_707 = core__GEN_9_1;
  assign _GEN_1455 = {_GEN_1454,profilePin_707}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_708 = core__GEN_10_2;
  assign _GEN_1456 = {_GEN_1455,profilePin_708}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_709 = core__GEN_11_1;
  assign _GEN_1457 = {_GEN_1456,profilePin_709}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_710 = core__GEN_12;
  assign _GEN_1458 = {_GEN_1457,profilePin_710}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_711 = core__GEN_13_0;
  assign _GEN_1459 = {_GEN_1458,profilePin_711}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_712 = core__GEN_14_0;
  assign _GEN_1460 = {_GEN_1459,profilePin_712}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_713 = core__GEN_15;
  assign _GEN_1461 = {_GEN_1460,profilePin_713}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_714 = core__GEN_16;
  assign _GEN_1462 = {_GEN_1461,profilePin_714}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_715 = core__GEN_17;
  assign _GEN_1463 = {_GEN_1462,profilePin_715}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_716 = core__GEN_18_0;
  assign _GEN_1464 = {_GEN_1463,profilePin_716}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_717 = core__GEN_19;
  assign _GEN_1465 = {_GEN_1464,profilePin_717}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_718 = core__GEN_20;
  assign _GEN_1466 = {_GEN_1465,profilePin_718}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_719 = core__GEN_21;
  assign _GEN_1467 = {_GEN_1466,profilePin_719}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_720 = core__GEN_22;
  assign _GEN_1468 = {_GEN_1467,profilePin_720}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_721 = core__GEN_23;
  assign _GEN_1469 = {_GEN_1468,profilePin_721}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_722 = memory__GEN_0_4;
  assign _GEN_1470 = {_GEN_1469,profilePin_722}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_723 = memory__GEN_1_3;
  assign _GEN_1471 = {_GEN_1470,profilePin_723}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_724 = memory__GEN_2_2;
  assign _GEN_1472 = {_GEN_1471,profilePin_724}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_725 = memory__GEN_3_0;
  assign _GEN_1473 = {_GEN_1472,profilePin_725}; // @[:Sodor3Stage.fir@3963.2]
  assign _GEN_1474 = {_GEN_1473,1'h1}; // @[:Sodor3Stage.fir@3963.2]
  assign _GEN_1475 = {_GEN_1474,1'h1}; // @[:Sodor3Stage.fir@3963.2]
  assign _GEN_1476 = {_GEN_1475,1'h1}; // @[:Sodor3Stage.fir@3963.2]
  assign _GEN_1477 = {_GEN_1476,1'h1}; // @[:Sodor3Stage.fir@3963.2]
  assign _GEN_1478 = {_GEN_1477,1'h1}; // @[:Sodor3Stage.fir@3963.2]
  assign _GEN_1479 = {_GEN_1478,1'h1}; // @[:Sodor3Stage.fir@3963.2]
  assign _GEN_1480 = {_GEN_1479,1'h1}; // @[:Sodor3Stage.fir@3963.2]
  assign _GEN_1481 = {_GEN_1480,1'h1}; // @[:Sodor3Stage.fir@3963.2]
  assign _GEN_1482 = {_GEN_1481,1'h1}; // @[:Sodor3Stage.fir@3963.2]
  assign _GEN_1483 = {_GEN_1482,1'h1}; // @[:Sodor3Stage.fir@3963.2]
  assign _GEN_1484 = {_GEN_1483,1'h1}; // @[:Sodor3Stage.fir@3963.2]
  assign _GEN_1485 = {_GEN_1484,1'h1}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_738 = memory__GEN_0_2;
  assign _GEN_1486 = {_GEN_1485,profilePin_738}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_739 = memory__GEN_1_1;
  assign _GEN_1487 = {_GEN_1486,profilePin_739}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_740 = memory__GEN_2_4;
  assign _GEN_1488 = {_GEN_1487,profilePin_740}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_741 = memory__GEN_3_4;
  assign _GEN_1489 = {_GEN_1488,profilePin_741}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_742 = memory__GEN_4_0;
  assign _GEN_1490 = {_GEN_1489,profilePin_742}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_743 = memory__GEN_5_6;
  assign _GEN_1491 = {_GEN_1490,profilePin_743}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_744 = memory__GEN_6_3;
  assign _GEN_1492 = {_GEN_1491,profilePin_744}; // @[:Sodor3Stage.fir@3963.2]
  assign profilePin_745 = memory__GEN_7_0;
  assign io_imem_req_valid = 1'h1;
  assign io_imem_req_bits_addr = core_io_imem_req_bits_addr;
  assign io_imem_req_bits_data = 32'h0;
  assign io_imem_req_bits_fcn = 1'h0;
  assign io_imem_req_bits_typ = 3'h7;
  assign assert_out = core__GEN_388;
  assign auto_cover_out = {_GEN_1492,profilePin_745};
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_imem_resp_bits_data = io_imem_resp_bits_data;
  assign core_io_dmem_resp_bits_data = memory_io_core_ports_0_resp_bits_data;
  assign memory_clock = clock;
  assign memory_io_core_ports_0_req_bits_addr = core_io_dmem_req_bits_addr;
  assign memory_io_core_ports_0_req_bits_data = core_io_dmem_req_bits_data;
  assign memory_io_core_ports_0_req_bits_fcn = core_io_dmem_req_bits_fcn;
  assign memory_io_core_ports_0_req_bits_typ = core_io_dmem_req_bits_typ;
endmodule
module FrontEnd( // @[:Sodor3Stage.fir@414.2]
  input         metaReset,
  input         clock, // @[:Sodor3Stage.fir@415.4]
  input         reset, // @[:Sodor3Stage.fir@416.4]
  input         io_cpu_req_valid, // @[:Sodor3Stage.fir@417.4]
  input  [31:0] io_cpu_req_bits_pc, // @[:Sodor3Stage.fir@417.4]
  input         io_cpu_resp_ready, // @[:Sodor3Stage.fir@417.4]
  output        io_cpu_resp_valid, // @[:Sodor3Stage.fir@417.4]
  output [31:0] io_cpu_resp_bits_pc, // @[:Sodor3Stage.fir@417.4]
  output [31:0] io_cpu_resp_bits_inst, // @[:Sodor3Stage.fir@417.4]
  output [31:0] io_imem_req_bits_addr, // @[:Sodor3Stage.fir@417.4]
  input  [31:0] io_imem_resp_bits_data, // @[:Sodor3Stage.fir@417.4]
  output        _GEN_1_0,
  output        _GEN_10_0,
  output        _GEN_13_0,
  output        _GEN_7_1,
  output        _GEN_9_4,
  output        _GEN_12_2,
  output        _GEN_6_4,
  output        _GEN_14_3,
  output        _GEN_5_4,
  output        _GEN_8_4,
  output        _GEN_11_4
);
  reg  if_reg_valid; // @[frontend.scala 87:27:Sodor3Stage.fir@435.4]
  reg [31:0] _RAND_0;
  reg [31:0] if_reg_pc; // @[frontend.scala 88:27:Sodor3Stage.fir@439.4]
  reg [31:0] _RAND_1;
  reg  exe_reg_valid; // @[frontend.scala 90:27:Sodor3Stage.fir@440.4]
  reg [31:0] _RAND_2;
  reg [31:0] exe_reg_pc; // @[frontend.scala 91:27:Sodor3Stage.fir@441.4]
  reg [31:0] _RAND_3;
  reg [31:0] exe_reg_inst; // @[frontend.scala 92:27:Sodor3Stage.fir@442.4]
  reg [31:0] _RAND_4;
  wire [32:0] _T_130; // @[frontend.scala 88:45:Sodor3Stage.fir@436.4]
  wire [32:0] _T_131; // @[frontend.scala 88:45:Sodor3Stage.fir@437.4]
  wire [31:0] _T_132; // @[frontend.scala 88:45:Sodor3Stage.fir@438.4]
  wire [32:0] _T_142; // @[frontend.scala 100:33:Sodor3Stage.fir@446.4]
  wire [31:0] if_pc_plus4; // @[frontend.scala 100:33:Sodor3Stage.fir@447.4]
  wire [31:0] _GEN_0; // @[frontend.scala 107:7:Sodor3Stage.fir@450.6]
  wire  _T_144; // @[frontend.scala 133:40:Sodor3Stage.fir@466.6]
  wire  _T_145; // @[frontend.scala 133:37:Sodor3Stage.fir@467.6]
  assign _T_130 = 32'h80000000 - 32'h4; // @[frontend.scala 88:45:Sodor3Stage.fir@436.4]
  assign _T_131 = $unsigned(_T_130); // @[frontend.scala 88:45:Sodor3Stage.fir@437.4]
  assign _T_132 = _T_131[31:0]; // @[frontend.scala 88:45:Sodor3Stage.fir@438.4]
  assign _T_142 = if_reg_pc + 32'h4; // @[frontend.scala 100:33:Sodor3Stage.fir@446.4]
  assign if_pc_plus4 = _T_142[31:0]; // @[frontend.scala 100:33:Sodor3Stage.fir@447.4]
  assign _GEN_0 = io_cpu_req_valid ? io_cpu_req_bits_pc : if_pc_plus4; // @[frontend.scala 107:7:Sodor3Stage.fir@450.6]
  assign _T_144 = io_cpu_req_valid == 1'h0; // @[frontend.scala 133:40:Sodor3Stage.fir@466.6]
  assign _T_145 = if_reg_valid & _T_144; // @[frontend.scala 133:37:Sodor3Stage.fir@467.6]
  assign io_cpu_resp_valid = exe_reg_valid;
  assign io_cpu_resp_bits_pc = exe_reg_pc;
  assign io_cpu_resp_bits_inst = exe_reg_inst;
  assign io_imem_req_bits_addr = io_cpu_resp_ready ? _GEN_0 : if_reg_pc;
  assign _GEN_1_0 = io_cpu_req_valid;
  assign _GEN_10_0 = reset;
  assign _GEN_13_0 = io_cpu_resp_ready;
  assign _GEN_7_1 = io_cpu_resp_ready;
  assign _GEN_9_4 = io_cpu_resp_ready;
  assign _GEN_12_2 = reset;
  assign _GEN_6_4 = io_cpu_resp_ready;
  assign _GEN_14_3 = io_cpu_resp_ready;
  assign _GEN_5_4 = io_cpu_resp_ready;
  assign _GEN_8_4 = io_cpu_resp_ready;
  assign _GEN_11_4 = reset;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  if_reg_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  if_reg_pc = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  exe_reg_valid = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  exe_reg_pc = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  exe_reg_inst = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (metaReset) begin
      if_reg_valid <= 1'h0;
    end else begin
      if (reset) begin
        if_reg_valid <= 1'h0;
      end else begin
        if (io_cpu_resp_ready) begin
          if_reg_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      if_reg_pc <= 32'h0;
    end else begin
      if (reset) begin
        if_reg_pc <= _T_132;
      end else begin
        if (io_cpu_resp_ready) begin
          if (io_cpu_resp_ready) begin
            if (io_cpu_req_valid) begin
              if_reg_pc <= io_cpu_req_bits_pc;
            end else begin
              if_reg_pc <= if_pc_plus4;
            end
          end
        end
      end
    end
    if (metaReset) begin
      exe_reg_valid <= 1'h0;
    end else begin
      if (reset) begin
        exe_reg_valid <= 1'h0;
      end else begin
        if (io_cpu_resp_ready) begin
          exe_reg_valid <= _T_145;
        end
      end
    end
    if (metaReset) begin
      exe_reg_pc <= 32'h0;
    end else begin
      if (io_cpu_resp_ready) begin
        exe_reg_pc <= if_reg_pc;
      end
    end
    if (metaReset) begin
      exe_reg_inst <= 32'h0;
    end else begin
      if (io_cpu_resp_ready) begin
        exe_reg_inst <= io_imem_resp_bits_data;
      end
    end
  end
endmodule
module CtlPath( // @[:Sodor3Stage.fir@478.2]
  input         metaReset,
  input         clock, // @[:Sodor3Stage.fir@479.4]
  output        io_imem_req_valid, // @[:Sodor3Stage.fir@481.4]
  input         io_imem_resp_valid, // @[:Sodor3Stage.fir@481.4]
  input  [31:0] io_imem_resp_bits_inst, // @[:Sodor3Stage.fir@481.4]
  input         io_dat_br_eq, // @[:Sodor3Stage.fir@481.4]
  input         io_dat_br_lt, // @[:Sodor3Stage.fir@481.4]
  input         io_dat_br_ltu, // @[:Sodor3Stage.fir@481.4]
  input         io_dat_csr_eret, // @[:Sodor3Stage.fir@481.4]
  output        io_ctl_exe_kill, // @[:Sodor3Stage.fir@481.4]
  output [2:0]  io_ctl_pc_sel, // @[:Sodor3Stage.fir@481.4]
  output        io_ctl_brjmp_sel, // @[:Sodor3Stage.fir@481.4]
  output [1:0]  io_ctl_op1_sel, // @[:Sodor3Stage.fir@481.4]
  output [1:0]  io_ctl_op2_sel, // @[:Sodor3Stage.fir@481.4]
  output [3:0]  io_ctl_alu_fun, // @[:Sodor3Stage.fir@481.4]
  output [1:0]  io_ctl_wb_sel, // @[:Sodor3Stage.fir@481.4]
  output        io_ctl_rf_wen, // @[:Sodor3Stage.fir@481.4]
  output        io_ctl_bypassable, // @[:Sodor3Stage.fir@481.4]
  output [2:0]  io_ctl_csr_cmd, // @[:Sodor3Stage.fir@481.4]
  output        io_ctl_dmem_fcn, // @[:Sodor3Stage.fir@481.4]
  output [2:0]  io_ctl_dmem_typ, // @[:Sodor3Stage.fir@481.4]
  output        io_ctl_exception, // @[:Sodor3Stage.fir@481.4]
  output        _GEN_91_0,
  output        _GEN_51_0,
  output        _GEN_304_0,
  output        _GEN_199_0,
  output        _GEN_148_0,
  output        _GEN_403_0,
  output        _GEN_24_0,
  output        _GEN_247_0,
  output        _GEN_106_0,
  output        _GEN_133_0,
  output        _GEN_205_0,
  output        _GEN_39_0,
  output        _GEN_232_0,
  output        _GEN_418_0,
  output        _GEN_127_0,
  output        _GEN_331_0,
  output        _GEN_190_0,
  output        _GEN_226_0,
  output        _GEN_45_0,
  output        _GEN_112_0,
  output        _GEN_298_0,
  output        _GEN_72_0,
  output        _GEN_211_0,
  output        _GEN_325_0,
  output        _GEN_397_0,
  output        _GEN_424_0,
  output        _GEN_30_0,
  output        _GEN_310_0,
  output        _GEN_319_0,
  output        _GEN_66_0,
  output        _GEN_220_0,
  output        _GEN_214_0,
  output        _GEN_100_0,
  output        _GEN_109_0,
  output        _GEN_313_0,
  output        _GEN_282_0,
  output        _GEN_177_0,
  output        _GEN_208_0,
  output        _GEN_391_0,
  output        _GEN_381_0,
  output        _GEN_412_0,
  output        _GEN_27_0,
  output        _GEN_276_0,
  output        _GEN_54_0,
  output        _GEN_193_0,
  output        _GEN_12_1,
  output        _GEN_406_0,
  output        _GEN_48_0,
  output        _GEN_115_0,
  output        _GEN_6_1,
  output        _GEN_33_0,
  output        _GEN_121_0,
  output        _GEN_307_0,
  output        _GEN_375_0,
  output        _GEN_229_0,
  output        _GEN_94_0,
  output        _GEN_292_0,
  output        _GEN_183_0,
  output        _GEN_0_1,
  output        _GEN_196_0,
  output        _GEN_186_0,
  output        _GEN_400_0,
  output        _GEN_103_0,
  output        _GEN_264_0,
  output        _GEN_295_0,
  output        _GEN_159_0,
  output        _GEN_202_0,
  output        _GEN_171_0,
  output        _GEN_357_0,
  output        _GEN_270_0,
  output        _GEN_384_0,
  output        _GEN_36_0,
  output        _GEN_285_0,
  output        _GEN_165_0,
  output        _GEN_279_0,
  output        _GEN_378_0,
  output        _GEN_21_1,
  output        _GEN_301_0,
  output        _GEN_394_0,
  output        _GEN_15_1,
  output        _GEN_363_0,
  output        _GEN_9_3,
  output        _GEN_258_0,
  output        _GEN_97_0,
  output        _GEN_345_0,
  output        _GEN_339_0,
  output        _GEN_18_0,
  output        _GEN_147_0,
  output        _GEN_330_0,
  output        _GEN_86_0,
  output        _GEN_273_0,
  output        _GEN_351_0,
  output        _GEN_231_0,
  output        _GEN_189_0,
  output        _GEN_153_0,
  output        _GEN_288_0,
  output        _GEN_366_0,
  output        _GEN_252_0,
  output        _GEN_180_0,
  output        _GEN_71_0,
  output        _GEN_174_0,
  output        _GEN_168_0,
  output        _GEN_372_0,
  output        _GEN_3_2,
  output        _GEN_387_0,
  output        _GEN_246_0,
  output        _GEN_267_0,
  output        _GEN_354_0,
  output        _GEN_213_0,
  output        _GEN_249_0,
  output        _GEN_240_0,
  output        _GEN_141_0,
  output        _GEN_135_0,
  output        _GEN_234_0,
  output        _GEN_348_0,
  output        _GEN_261_0,
  output        _GEN_312_0,
  output        _GEN_53_0,
  output        _GEN_333_0,
  output        _GEN_68_0,
  output        _GEN_156_0,
  output        _GEN_360_0,
  output        _GEN_369_0,
  output        _GEN_74_0,
  output        _GEN_327_0,
  output        _GEN_89_0,
  output        _GEN_162_0,
  output        _GEN_426_0,
  output        _GEN_129_0,
  output        _GEN_228_0,
  output        _GEN_411_0,
  output        _GEN_255_0,
  output        _GEN_120_0,
  output        _GEN_80_0,
  output        _GEN_342_0,
  output        _GEN_393_0,
  output        _GEN_56_0,
  output        _GEN_144_0,
  output        _GEN_408_0,
  output        _GEN_222_0,
  output        _GEN_117_0,
  output        _GEN_321_0,
  output        _GEN_243_0,
  output        _GEN_237_0,
  output        _GEN_123_0,
  output        _GEN_102_0,
  output        _GEN_62_0,
  output        _GEN_150_0,
  output        _GEN_336_0,
  output        _GEN_201_0,
  output        _GEN_195_0,
  output        _GEN_414_0,
  output        _GEN_300_0,
  output        _GEN_294_0,
  output        _GEN_309_0,
  output        _GEN_77_0,
  output        _GEN_83_0,
  output        _GEN_216_0,
  output        _GEN_420_0,
  output        _GEN_35_0,
  output        _GEN_41_0,
  output        _GEN_315_0,
  output        _GEN_429_0,
  output        _GEN_138_0,
  output        _GEN_402_0,
  output        _GEN_17_1,
  output        _GEN_225_0,
  output        _GEN_105_0,
  output        _GEN_50_0,
  output        _GEN_44_0,
  output        _GEN_324_0,
  output        _GEN_318_0,
  output        _GEN_396_0,
  output        _GEN_386_0,
  output        _GEN_38_0,
  output        _GEN_65_0,
  output        _GEN_23_1,
  output        _GEN_417_0,
  output        _GEN_111_0,
  output        _GEN_210_0,
  output        _GEN_219_0,
  output        _GEN_423_0,
  output        _GEN_132_0,
  output        _GEN_126_0,
  output        _GEN_287_0,
  output        _GEN_90_0,
  output        _GEN_204_0,
  output        _GEN_99_0,
  output        _GEN_303_0,
  output        _GEN_297_0,
  output        _GEN_59_0,
  output        _GEN_188_0,
  output        _GEN_198_0,
  output        _GEN_176_0,
  output        _GEN_11_3,
  output        _GEN_380_0,
  output        _GEN_93_0,
  output        _GEN_161_0,
  output        _GEN_192_0,
  output        _GEN_207_0,
  output        _GEN_405_0,
  output        _GEN_260_0,
  output        _GEN_26_0,
  output        _GEN_114_0,
  output        _GEN_269_0,
  output        _GEN_182_0,
  output        _GEN_399_0,
  output        _GEN_368_0,
  output        _GEN_390_0,
  output        _GEN_32_0,
  output        _GEN_281_0,
  output        _GEN_275_0,
  output        _GEN_291_0,
  output        _GEN_47_0,
  output        _GEN_5_3,
  output        _GEN_389_0,
  output        _GEN_306_0,
  output        _GEN_374_0,
  output        _GEN_108_0,
  output        _GEN_356_0,
  output        _GEN_20_1,
  output        _GEN_14_2,
  output        _GEN_29_0,
  output        _GEN_82_0,
  output        _GEN_170_0,
  output        _GEN_185_0,
  output        _GEN_278_0,
  output        _GEN_143_0,
  output        _GEN_96_0,
  output        _GEN_263_0,
  output        _GEN_164_0,
  output        _GEN_158_0,
  output        _GEN_362_0,
  output        _GEN_377_0,
  output        _GEN_257_0,
  output        _GEN_284_0,
  output        _GEN_179_0,
  output        _GEN_383_0,
  output        _GEN_242_0,
  output        _GEN_8_3,
  output        _GEN_341_0,
  output        _GEN_76_0,
  output        _GEN_173_0,
  output        _GEN_224_1,
  output        _GEN_359_0,
  output        _GEN_251_0,
  output        _GEN_131_0,
  output        _GEN_146_0,
  output        _GEN_350_0,
  output        _GEN_344_0,
  output        _GEN_239_1,
  output        _GEN_272_0,
  output        _GEN_64_0,
  output        _GEN_58_0,
  output        _GEN_230_0,
  output        _GEN_365_0,
  output        _GEN_323_1,
  output        _GEN_85_0,
  output        _GEN_338_1,
  output        _GEN_79_0,
  output        _GEN_2_3,
  output        _GEN_245_0,
  output        _GEN_70_0,
  output        _GEN_152_0,
  output        _GEN_167_0,
  output        _GEN_422_0,
  output        _GEN_371_0,
  output        _GEN_266_0,
  output        _GEN_125_0,
  output        _GEN_212_1,
  output        _GEN_254_0,
  output        _GEN_155_0,
  output        _GEN_149_0,
  output        _GEN_227_0,
  output        _GEN_113_0,
  output        _GEN_140_0,
  output        _GEN_326_0,
  output        _GEN_425_0,
  output        _GEN_404_0,
  output        _GEN_353_0,
  output        _GEN_248_0,
  output        _GEN_107_0,
  output        _GEN_311_1,
  output        _GEN_73_0,
  output        _GEN_67_0,
  output        _GEN_347_0,
  output        _GEN_206_1,
  output        _GEN_410_0,
  output        _GEN_419_0,
  output        _GEN_233_0,
  output        _GEN_305_1,
  output        _GEN_128_0,
  output        _GEN_332_0,
  output        _GEN_88_0,
  output        _GEN_52_0,
  output        _GEN_46_0,
  output        _GEN_134_0,
  output        _GEN_221_0,
  output        _GEN_407_0,
  output        _GEN_382_1,
  output        _GEN_28_0,
  output        _GEN_40_0,
  output        _GEN_55_0,
  output        _GEN_329_0,
  output        _GEN_194_1,
  output        _GEN_392_0,
  output        _GEN_236_0,
  output        _GEN_101_0,
  output        _GEN_61_0,
  output        _GEN_34_0,
  output        _GEN_116_0,
  output        _GEN_122_0,
  output        _GEN_320_1,
  output        _GEN_215_0,
  output        _GEN_335_0,
  output        _GEN_293_1,
  output        _GEN_428_0,
  output        _GEN_49_0,
  output        _GEN_137_0,
  output        _GEN_200_1,
  output        _GEN_209_0,
  output        _GEN_95_0,
  output        _GEN_413_0,
  output        _GEN_314_0,
  output        _GEN_308_0,
  output        _GEN_16_1,
  output        _GEN_395_0,
  output        _GEN_385_1,
  output        _GEN_104_0,
  output        _GEN_302_1,
  output        _GEN_317_1,
  output        _GEN_203_1,
  output        _GEN_172_1,
  output        _GEN_197_1,
  output        _GEN_370_1,
  output        _GEN_416_0,
  output        _GEN_22_1,
  output        _GEN_271_1,
  output        _GEN_119_0,
  output        _GEN_379_1,
  output        _GEN_187_1,
  output        _GEN_401_0,
  output        _GEN_43_0,
  output        _GEN_296_1,
  output        _GEN_286_1,
  output        _GEN_364_1,
  output        _GEN_1_5,
  output        _GEN_98_0,
  output        _GEN_37_0,
  output        _GEN_110_0,
  output        _GEN_218_1,
  output        _GEN_25_0,
  output        _GEN_181_1,
  output        _GEN_175_1,
  output        _GEN_289_1,
  output        _GEN_352_1,
  output        _GEN_31_0,
  output        _GEN_274_1,
  output        _GEN_160_1,
  output        _GEN_169_1,
  output        _GEN_191_1,
  output        _GEN_373_1,
  output        _GEN_19_1,
  output        _GEN_367_1,
  output        _GEN_268_1,
  output        _GEN_290_1,
  output        _GEN_280_1,
  output        _GEN_154_1,
  output        _GEN_87_0,
  output        _GEN_299_1,
  output        _GEN_10_4,
  output        _GEN_398_0,
  output        _GEN_4_4,
  output        _GEN_388_1,
  output        _GEN_253_1,
  output        _GEN_92_0,
  output        _GEN_346_1,
  output        _GEN_334_1,
  output        _GEN_340_1,
  output        _GEN_13_3,
  output        _GEN_256_1,
  output        _GEN_328_1,
  output        _GEN_81_0,
  output        _GEN_355_1,
  output        _GEN_7_6,
  output        _GEN_277_1,
  output        _GEN_69_0,
  output        _GEN_157_1,
  output        _GEN_235_1,
  output        _GEN_184_1,
  output        _GEN_60_0,
  output        _GEN_283_1,
  output        _GEN_142_0,
  output        _GEN_178_1,
  output        _GEN_241_1,
  output        _GEN_361_1,
  output        _GEN_136_0,
  output        _GEN_75_0,
  output        _GEN_163_1,
  output        _GEN_349_1,
  output        _GEN_427_0,
  output        _GEN_376_1,
  output        _GEN_262_1,
  output        _GEN_166_1,
  output        _GEN_358_1,
  output        _GEN_42_0,
  output        _GEN_265_1,
  output        _GEN_316_1,
  output        _GEN_130_0,
  output        _GEN_124_0,
  output        _GEN_343_1,
  output        _GEN_223_1,
  output        _GEN_238_1,
  output        _GEN_118_0,
  output        _GEN_151_1,
  output        _GEN_145_0,
  output        _GEN_337_1,
  output        _GEN_244_1,
  output        _GEN_409_0,
  output        _GEN_322_1,
  output        _GEN_78_0,
  output        _GEN_217_1,
  output        _GEN_421_0,
  output        _GEN_415_0,
  output        _GEN_63_0,
  output        _GEN_57_0,
  output        _GEN_250_1,
  output        _GEN_259_1,
  output        _GEN_139_0,
  output        _GEN_84_0
);
  reg  _T_1028; // @[cpath.scala 179:27:Sodor3Stage.fir@1383.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@518.4]
  wire  _T_89; // @[Lookup.scala 9:38:Sodor3Stage.fir@519.4]
  wire  _T_93; // @[Lookup.scala 9:38:Sodor3Stage.fir@521.4]
  wire  _T_97; // @[Lookup.scala 9:38:Sodor3Stage.fir@523.4]
  wire  _T_101; // @[Lookup.scala 9:38:Sodor3Stage.fir@525.4]
  wire  _T_105; // @[Lookup.scala 9:38:Sodor3Stage.fir@527.4]
  wire  _T_109; // @[Lookup.scala 9:38:Sodor3Stage.fir@529.4]
  wire  _T_113; // @[Lookup.scala 9:38:Sodor3Stage.fir@531.4]
  wire  _T_117; // @[Lookup.scala 9:38:Sodor3Stage.fir@533.4]
  wire [31:0] _T_120; // @[Lookup.scala 9:38:Sodor3Stage.fir@534.4]
  wire  _T_121; // @[Lookup.scala 9:38:Sodor3Stage.fir@535.4]
  wire  _T_125; // @[Lookup.scala 9:38:Sodor3Stage.fir@537.4]
  wire  _T_129; // @[Lookup.scala 9:38:Sodor3Stage.fir@539.4]
  wire  _T_133; // @[Lookup.scala 9:38:Sodor3Stage.fir@541.4]
  wire  _T_137; // @[Lookup.scala 9:38:Sodor3Stage.fir@543.4]
  wire  _T_141; // @[Lookup.scala 9:38:Sodor3Stage.fir@545.4]
  wire  _T_145; // @[Lookup.scala 9:38:Sodor3Stage.fir@547.4]
  wire  _T_149; // @[Lookup.scala 9:38:Sodor3Stage.fir@549.4]
  wire [31:0] _T_152; // @[Lookup.scala 9:38:Sodor3Stage.fir@550.4]
  wire  _T_153; // @[Lookup.scala 9:38:Sodor3Stage.fir@551.4]
  wire  _T_157; // @[Lookup.scala 9:38:Sodor3Stage.fir@553.4]
  wire  _T_161; // @[Lookup.scala 9:38:Sodor3Stage.fir@555.4]
  wire [31:0] _T_164; // @[Lookup.scala 9:38:Sodor3Stage.fir@556.4]
  wire  _T_165; // @[Lookup.scala 9:38:Sodor3Stage.fir@557.4]
  wire  _T_169; // @[Lookup.scala 9:38:Sodor3Stage.fir@559.4]
  wire  _T_173; // @[Lookup.scala 9:38:Sodor3Stage.fir@561.4]
  wire  _T_177; // @[Lookup.scala 9:38:Sodor3Stage.fir@563.4]
  wire  _T_181; // @[Lookup.scala 9:38:Sodor3Stage.fir@565.4]
  wire  _T_185; // @[Lookup.scala 9:38:Sodor3Stage.fir@567.4]
  wire  _T_189; // @[Lookup.scala 9:38:Sodor3Stage.fir@569.4]
  wire  _T_193; // @[Lookup.scala 9:38:Sodor3Stage.fir@571.4]
  wire  _T_197; // @[Lookup.scala 9:38:Sodor3Stage.fir@573.4]
  wire  _T_201; // @[Lookup.scala 9:38:Sodor3Stage.fir@575.4]
  wire  _T_205; // @[Lookup.scala 9:38:Sodor3Stage.fir@577.4]
  wire  _T_209; // @[Lookup.scala 9:38:Sodor3Stage.fir@579.4]
  wire  _T_213; // @[Lookup.scala 9:38:Sodor3Stage.fir@581.4]
  wire  _T_217; // @[Lookup.scala 9:38:Sodor3Stage.fir@583.4]
  wire  _T_221; // @[Lookup.scala 9:38:Sodor3Stage.fir@585.4]
  wire  _T_225; // @[Lookup.scala 9:38:Sodor3Stage.fir@587.4]
  wire  _T_229; // @[Lookup.scala 9:38:Sodor3Stage.fir@589.4]
  wire  _T_233; // @[Lookup.scala 9:38:Sodor3Stage.fir@591.4]
  wire  _T_237; // @[Lookup.scala 9:38:Sodor3Stage.fir@593.4]
  wire  _T_241; // @[Lookup.scala 9:38:Sodor3Stage.fir@595.4]
  wire  _T_245; // @[Lookup.scala 9:38:Sodor3Stage.fir@597.4]
  wire  _T_249; // @[Lookup.scala 9:38:Sodor3Stage.fir@599.4]
  wire  _T_253; // @[Lookup.scala 9:38:Sodor3Stage.fir@601.4]
  wire  _T_257; // @[Lookup.scala 9:38:Sodor3Stage.fir@603.4]
  wire  _T_261; // @[Lookup.scala 9:38:Sodor3Stage.fir@605.4]
  wire  _T_265; // @[Lookup.scala 9:38:Sodor3Stage.fir@607.4]
  wire  _T_269; // @[Lookup.scala 9:38:Sodor3Stage.fir@609.4]
  wire  _T_273; // @[Lookup.scala 9:38:Sodor3Stage.fir@611.4]
  wire  _T_277; // @[Lookup.scala 9:38:Sodor3Stage.fir@613.4]
  wire  _T_281; // @[Lookup.scala 9:38:Sodor3Stage.fir@615.4]
  wire  _T_285; // @[Lookup.scala 9:38:Sodor3Stage.fir@617.4]
  wire  _T_287; // @[Lookup.scala 11:37:Sodor3Stage.fir@619.4]
  wire  _T_288; // @[Lookup.scala 11:37:Sodor3Stage.fir@620.4]
  wire  _T_289; // @[Lookup.scala 11:37:Sodor3Stage.fir@621.4]
  wire  _T_290; // @[Lookup.scala 11:37:Sodor3Stage.fir@622.4]
  wire  _T_291; // @[Lookup.scala 11:37:Sodor3Stage.fir@623.4]
  wire  _T_292; // @[Lookup.scala 11:37:Sodor3Stage.fir@624.4]
  wire  _T_293; // @[Lookup.scala 11:37:Sodor3Stage.fir@625.4]
  wire  _T_294; // @[Lookup.scala 11:37:Sodor3Stage.fir@626.4]
  wire  _T_295; // @[Lookup.scala 11:37:Sodor3Stage.fir@627.4]
  wire  _T_296; // @[Lookup.scala 11:37:Sodor3Stage.fir@628.4]
  wire  _T_297; // @[Lookup.scala 11:37:Sodor3Stage.fir@629.4]
  wire  _T_298; // @[Lookup.scala 11:37:Sodor3Stage.fir@630.4]
  wire  _T_299; // @[Lookup.scala 11:37:Sodor3Stage.fir@631.4]
  wire  _T_300; // @[Lookup.scala 11:37:Sodor3Stage.fir@632.4]
  wire  _T_301; // @[Lookup.scala 11:37:Sodor3Stage.fir@633.4]
  wire  _T_302; // @[Lookup.scala 11:37:Sodor3Stage.fir@634.4]
  wire  _T_303; // @[Lookup.scala 11:37:Sodor3Stage.fir@635.4]
  wire  _T_304; // @[Lookup.scala 11:37:Sodor3Stage.fir@636.4]
  wire  _T_305; // @[Lookup.scala 11:37:Sodor3Stage.fir@637.4]
  wire  _T_306; // @[Lookup.scala 11:37:Sodor3Stage.fir@638.4]
  wire  _T_307; // @[Lookup.scala 11:37:Sodor3Stage.fir@639.4]
  wire  _T_308; // @[Lookup.scala 11:37:Sodor3Stage.fir@640.4]
  wire  _T_309; // @[Lookup.scala 11:37:Sodor3Stage.fir@641.4]
  wire  _T_310; // @[Lookup.scala 11:37:Sodor3Stage.fir@642.4]
  wire  _T_311; // @[Lookup.scala 11:37:Sodor3Stage.fir@643.4]
  wire  _T_312; // @[Lookup.scala 11:37:Sodor3Stage.fir@644.4]
  wire  _T_313; // @[Lookup.scala 11:37:Sodor3Stage.fir@645.4]
  wire  _T_314; // @[Lookup.scala 11:37:Sodor3Stage.fir@646.4]
  wire  _T_315; // @[Lookup.scala 11:37:Sodor3Stage.fir@647.4]
  wire  _T_316; // @[Lookup.scala 11:37:Sodor3Stage.fir@648.4]
  wire  _T_317; // @[Lookup.scala 11:37:Sodor3Stage.fir@649.4]
  wire  _T_318; // @[Lookup.scala 11:37:Sodor3Stage.fir@650.4]
  wire  _T_319; // @[Lookup.scala 11:37:Sodor3Stage.fir@651.4]
  wire  _T_320; // @[Lookup.scala 11:37:Sodor3Stage.fir@652.4]
  wire  _T_321; // @[Lookup.scala 11:37:Sodor3Stage.fir@653.4]
  wire  _T_322; // @[Lookup.scala 11:37:Sodor3Stage.fir@654.4]
  wire  _T_323; // @[Lookup.scala 11:37:Sodor3Stage.fir@655.4]
  wire  _T_324; // @[Lookup.scala 11:37:Sodor3Stage.fir@656.4]
  wire  _T_325; // @[Lookup.scala 11:37:Sodor3Stage.fir@657.4]
  wire  _T_326; // @[Lookup.scala 11:37:Sodor3Stage.fir@658.4]
  wire  _T_327; // @[Lookup.scala 11:37:Sodor3Stage.fir@659.4]
  wire  _T_328; // @[Lookup.scala 11:37:Sodor3Stage.fir@660.4]
  wire  _T_329; // @[Lookup.scala 11:37:Sodor3Stage.fir@661.4]
  wire  _T_330; // @[Lookup.scala 11:37:Sodor3Stage.fir@662.4]
  wire  _T_331; // @[Lookup.scala 11:37:Sodor3Stage.fir@663.4]
  wire  _T_332; // @[Lookup.scala 11:37:Sodor3Stage.fir@664.4]
  wire  _T_333; // @[Lookup.scala 11:37:Sodor3Stage.fir@665.4]
  wire  _T_334; // @[Lookup.scala 11:37:Sodor3Stage.fir@666.4]
  wire  cs_inst_val; // @[Lookup.scala 11:37:Sodor3Stage.fir@667.4]
  wire [3:0] _T_348; // @[Lookup.scala 11:37:Sodor3Stage.fir@681.4]
  wire [3:0] _T_349; // @[Lookup.scala 11:37:Sodor3Stage.fir@682.4]
  wire [3:0] _T_350; // @[Lookup.scala 11:37:Sodor3Stage.fir@683.4]
  wire [3:0] _T_351; // @[Lookup.scala 11:37:Sodor3Stage.fir@684.4]
  wire [3:0] _T_352; // @[Lookup.scala 11:37:Sodor3Stage.fir@685.4]
  wire [3:0] _T_353; // @[Lookup.scala 11:37:Sodor3Stage.fir@686.4]
  wire [3:0] _T_354; // @[Lookup.scala 11:37:Sodor3Stage.fir@687.4]
  wire [3:0] _T_355; // @[Lookup.scala 11:37:Sodor3Stage.fir@688.4]
  wire [3:0] _T_356; // @[Lookup.scala 11:37:Sodor3Stage.fir@689.4]
  wire [3:0] _T_357; // @[Lookup.scala 11:37:Sodor3Stage.fir@690.4]
  wire [3:0] _T_358; // @[Lookup.scala 11:37:Sodor3Stage.fir@691.4]
  wire [3:0] _T_359; // @[Lookup.scala 11:37:Sodor3Stage.fir@692.4]
  wire [3:0] _T_360; // @[Lookup.scala 11:37:Sodor3Stage.fir@693.4]
  wire [3:0] _T_361; // @[Lookup.scala 11:37:Sodor3Stage.fir@694.4]
  wire [3:0] _T_362; // @[Lookup.scala 11:37:Sodor3Stage.fir@695.4]
  wire [3:0] _T_363; // @[Lookup.scala 11:37:Sodor3Stage.fir@696.4]
  wire [3:0] _T_364; // @[Lookup.scala 11:37:Sodor3Stage.fir@697.4]
  wire [3:0] _T_365; // @[Lookup.scala 11:37:Sodor3Stage.fir@698.4]
  wire [3:0] _T_366; // @[Lookup.scala 11:37:Sodor3Stage.fir@699.4]
  wire [3:0] _T_367; // @[Lookup.scala 11:37:Sodor3Stage.fir@700.4]
  wire [3:0] _T_368; // @[Lookup.scala 11:37:Sodor3Stage.fir@701.4]
  wire [3:0] _T_369; // @[Lookup.scala 11:37:Sodor3Stage.fir@702.4]
  wire [3:0] _T_370; // @[Lookup.scala 11:37:Sodor3Stage.fir@703.4]
  wire [3:0] _T_371; // @[Lookup.scala 11:37:Sodor3Stage.fir@704.4]
  wire [3:0] _T_372; // @[Lookup.scala 11:37:Sodor3Stage.fir@705.4]
  wire [3:0] _T_373; // @[Lookup.scala 11:37:Sodor3Stage.fir@706.4]
  wire [3:0] _T_374; // @[Lookup.scala 11:37:Sodor3Stage.fir@707.4]
  wire [3:0] _T_375; // @[Lookup.scala 11:37:Sodor3Stage.fir@708.4]
  wire [3:0] _T_376; // @[Lookup.scala 11:37:Sodor3Stage.fir@709.4]
  wire [3:0] _T_377; // @[Lookup.scala 11:37:Sodor3Stage.fir@710.4]
  wire [3:0] _T_378; // @[Lookup.scala 11:37:Sodor3Stage.fir@711.4]
  wire [3:0] _T_379; // @[Lookup.scala 11:37:Sodor3Stage.fir@712.4]
  wire [3:0] _T_380; // @[Lookup.scala 11:37:Sodor3Stage.fir@713.4]
  wire [3:0] _T_381; // @[Lookup.scala 11:37:Sodor3Stage.fir@714.4]
  wire [3:0] _T_382; // @[Lookup.scala 11:37:Sodor3Stage.fir@715.4]
  wire [3:0] _T_383; // @[Lookup.scala 11:37:Sodor3Stage.fir@716.4]
  wire [3:0] cs_br_type; // @[Lookup.scala 11:37:Sodor3Stage.fir@717.4]
  wire  _T_404; // @[Lookup.scala 11:37:Sodor3Stage.fir@738.4]
  wire  _T_405; // @[Lookup.scala 11:37:Sodor3Stage.fir@739.4]
  wire  _T_406; // @[Lookup.scala 11:37:Sodor3Stage.fir@740.4]
  wire  _T_407; // @[Lookup.scala 11:37:Sodor3Stage.fir@741.4]
  wire  _T_408; // @[Lookup.scala 11:37:Sodor3Stage.fir@742.4]
  wire  _T_409; // @[Lookup.scala 11:37:Sodor3Stage.fir@743.4]
  wire  _T_410; // @[Lookup.scala 11:37:Sodor3Stage.fir@744.4]
  wire  _T_411; // @[Lookup.scala 11:37:Sodor3Stage.fir@745.4]
  wire  _T_412; // @[Lookup.scala 11:37:Sodor3Stage.fir@746.4]
  wire  _T_413; // @[Lookup.scala 11:37:Sodor3Stage.fir@747.4]
  wire  _T_414; // @[Lookup.scala 11:37:Sodor3Stage.fir@748.4]
  wire  _T_415; // @[Lookup.scala 11:37:Sodor3Stage.fir@749.4]
  wire  _T_416; // @[Lookup.scala 11:37:Sodor3Stage.fir@750.4]
  wire  _T_417; // @[Lookup.scala 11:37:Sodor3Stage.fir@751.4]
  wire  _T_418; // @[Lookup.scala 11:37:Sodor3Stage.fir@752.4]
  wire  _T_419; // @[Lookup.scala 11:37:Sodor3Stage.fir@753.4]
  wire  _T_420; // @[Lookup.scala 11:37:Sodor3Stage.fir@754.4]
  wire  _T_421; // @[Lookup.scala 11:37:Sodor3Stage.fir@755.4]
  wire  _T_422; // @[Lookup.scala 11:37:Sodor3Stage.fir@756.4]
  wire  _T_423; // @[Lookup.scala 11:37:Sodor3Stage.fir@757.4]
  wire  _T_424; // @[Lookup.scala 11:37:Sodor3Stage.fir@758.4]
  wire  _T_425; // @[Lookup.scala 11:37:Sodor3Stage.fir@759.4]
  wire  _T_426; // @[Lookup.scala 11:37:Sodor3Stage.fir@760.4]
  wire  _T_427; // @[Lookup.scala 11:37:Sodor3Stage.fir@761.4]
  wire  _T_428; // @[Lookup.scala 11:37:Sodor3Stage.fir@762.4]
  wire  _T_429; // @[Lookup.scala 11:37:Sodor3Stage.fir@763.4]
  wire  _T_430; // @[Lookup.scala 11:37:Sodor3Stage.fir@764.4]
  wire  _T_431; // @[Lookup.scala 11:37:Sodor3Stage.fir@765.4]
  wire  _T_432; // @[Lookup.scala 11:37:Sodor3Stage.fir@766.4]
  wire [1:0] _T_440; // @[Lookup.scala 11:37:Sodor3Stage.fir@775.4]
  wire [1:0] _T_441; // @[Lookup.scala 11:37:Sodor3Stage.fir@776.4]
  wire [1:0] _T_442; // @[Lookup.scala 11:37:Sodor3Stage.fir@777.4]
  wire [1:0] _T_443; // @[Lookup.scala 11:37:Sodor3Stage.fir@778.4]
  wire [1:0] _T_444; // @[Lookup.scala 11:37:Sodor3Stage.fir@779.4]
  wire [1:0] _T_445; // @[Lookup.scala 11:37:Sodor3Stage.fir@780.4]
  wire [1:0] _T_446; // @[Lookup.scala 11:37:Sodor3Stage.fir@781.4]
  wire [1:0] _T_447; // @[Lookup.scala 11:37:Sodor3Stage.fir@782.4]
  wire [1:0] _T_448; // @[Lookup.scala 11:37:Sodor3Stage.fir@783.4]
  wire [1:0] _T_449; // @[Lookup.scala 11:37:Sodor3Stage.fir@784.4]
  wire [1:0] _T_450; // @[Lookup.scala 11:37:Sodor3Stage.fir@785.4]
  wire [1:0] _T_451; // @[Lookup.scala 11:37:Sodor3Stage.fir@786.4]
  wire [1:0] _T_452; // @[Lookup.scala 11:37:Sodor3Stage.fir@787.4]
  wire [1:0] _T_453; // @[Lookup.scala 11:37:Sodor3Stage.fir@788.4]
  wire [1:0] _T_454; // @[Lookup.scala 11:37:Sodor3Stage.fir@789.4]
  wire [1:0] _T_455; // @[Lookup.scala 11:37:Sodor3Stage.fir@790.4]
  wire [1:0] _T_456; // @[Lookup.scala 11:37:Sodor3Stage.fir@791.4]
  wire [1:0] _T_457; // @[Lookup.scala 11:37:Sodor3Stage.fir@792.4]
  wire [1:0] _T_458; // @[Lookup.scala 11:37:Sodor3Stage.fir@793.4]
  wire [1:0] _T_459; // @[Lookup.scala 11:37:Sodor3Stage.fir@794.4]
  wire [1:0] _T_460; // @[Lookup.scala 11:37:Sodor3Stage.fir@795.4]
  wire [1:0] _T_461; // @[Lookup.scala 11:37:Sodor3Stage.fir@796.4]
  wire [1:0] _T_462; // @[Lookup.scala 11:37:Sodor3Stage.fir@797.4]
  wire [1:0] _T_463; // @[Lookup.scala 11:37:Sodor3Stage.fir@798.4]
  wire [1:0] _T_464; // @[Lookup.scala 11:37:Sodor3Stage.fir@799.4]
  wire [1:0] _T_465; // @[Lookup.scala 11:37:Sodor3Stage.fir@800.4]
  wire [1:0] _T_466; // @[Lookup.scala 11:37:Sodor3Stage.fir@801.4]
  wire [1:0] _T_467; // @[Lookup.scala 11:37:Sodor3Stage.fir@802.4]
  wire [1:0] _T_468; // @[Lookup.scala 11:37:Sodor3Stage.fir@803.4]
  wire [1:0] _T_469; // @[Lookup.scala 11:37:Sodor3Stage.fir@804.4]
  wire [1:0] _T_470; // @[Lookup.scala 11:37:Sodor3Stage.fir@805.4]
  wire [1:0] _T_471; // @[Lookup.scala 11:37:Sodor3Stage.fir@806.4]
  wire [1:0] _T_472; // @[Lookup.scala 11:37:Sodor3Stage.fir@807.4]
  wire [1:0] _T_473; // @[Lookup.scala 11:37:Sodor3Stage.fir@808.4]
  wire [1:0] _T_474; // @[Lookup.scala 11:37:Sodor3Stage.fir@809.4]
  wire [1:0] _T_475; // @[Lookup.scala 11:37:Sodor3Stage.fir@810.4]
  wire [1:0] _T_476; // @[Lookup.scala 11:37:Sodor3Stage.fir@811.4]
  wire [1:0] _T_477; // @[Lookup.scala 11:37:Sodor3Stage.fir@812.4]
  wire [1:0] _T_478; // @[Lookup.scala 11:37:Sodor3Stage.fir@813.4]
  wire [1:0] _T_479; // @[Lookup.scala 11:37:Sodor3Stage.fir@814.4]
  wire [1:0] _T_480; // @[Lookup.scala 11:37:Sodor3Stage.fir@815.4]
  wire [1:0] _T_481; // @[Lookup.scala 11:37:Sodor3Stage.fir@816.4]
  wire [1:0] _T_501; // @[Lookup.scala 11:37:Sodor3Stage.fir@837.4]
  wire [1:0] _T_502; // @[Lookup.scala 11:37:Sodor3Stage.fir@838.4]
  wire [1:0] _T_503; // @[Lookup.scala 11:37:Sodor3Stage.fir@839.4]
  wire [1:0] _T_504; // @[Lookup.scala 11:37:Sodor3Stage.fir@840.4]
  wire [1:0] _T_505; // @[Lookup.scala 11:37:Sodor3Stage.fir@841.4]
  wire [1:0] _T_506; // @[Lookup.scala 11:37:Sodor3Stage.fir@842.4]
  wire [1:0] _T_507; // @[Lookup.scala 11:37:Sodor3Stage.fir@843.4]
  wire [1:0] _T_508; // @[Lookup.scala 11:37:Sodor3Stage.fir@844.4]
  wire [1:0] _T_509; // @[Lookup.scala 11:37:Sodor3Stage.fir@845.4]
  wire [1:0] _T_510; // @[Lookup.scala 11:37:Sodor3Stage.fir@846.4]
  wire [1:0] _T_511; // @[Lookup.scala 11:37:Sodor3Stage.fir@847.4]
  wire [1:0] _T_512; // @[Lookup.scala 11:37:Sodor3Stage.fir@848.4]
  wire [1:0] _T_513; // @[Lookup.scala 11:37:Sodor3Stage.fir@849.4]
  wire [1:0] _T_514; // @[Lookup.scala 11:37:Sodor3Stage.fir@850.4]
  wire [1:0] _T_515; // @[Lookup.scala 11:37:Sodor3Stage.fir@851.4]
  wire [1:0] _T_516; // @[Lookup.scala 11:37:Sodor3Stage.fir@852.4]
  wire [1:0] _T_517; // @[Lookup.scala 11:37:Sodor3Stage.fir@853.4]
  wire [1:0] _T_518; // @[Lookup.scala 11:37:Sodor3Stage.fir@854.4]
  wire [1:0] _T_519; // @[Lookup.scala 11:37:Sodor3Stage.fir@855.4]
  wire [1:0] _T_520; // @[Lookup.scala 11:37:Sodor3Stage.fir@856.4]
  wire [1:0] _T_521; // @[Lookup.scala 11:37:Sodor3Stage.fir@857.4]
  wire [1:0] _T_522; // @[Lookup.scala 11:37:Sodor3Stage.fir@858.4]
  wire [1:0] _T_523; // @[Lookup.scala 11:37:Sodor3Stage.fir@859.4]
  wire [1:0] _T_524; // @[Lookup.scala 11:37:Sodor3Stage.fir@860.4]
  wire [1:0] _T_525; // @[Lookup.scala 11:37:Sodor3Stage.fir@861.4]
  wire [1:0] _T_526; // @[Lookup.scala 11:37:Sodor3Stage.fir@862.4]
  wire [1:0] _T_527; // @[Lookup.scala 11:37:Sodor3Stage.fir@863.4]
  wire [1:0] _T_528; // @[Lookup.scala 11:37:Sodor3Stage.fir@864.4]
  wire [1:0] _T_529; // @[Lookup.scala 11:37:Sodor3Stage.fir@865.4]
  wire [1:0] _T_530; // @[Lookup.scala 11:37:Sodor3Stage.fir@866.4]
  wire [3:0] _T_538; // @[Lookup.scala 11:37:Sodor3Stage.fir@875.4]
  wire [3:0] _T_539; // @[Lookup.scala 11:37:Sodor3Stage.fir@876.4]
  wire [3:0] _T_540; // @[Lookup.scala 11:37:Sodor3Stage.fir@877.4]
  wire [3:0] _T_541; // @[Lookup.scala 11:37:Sodor3Stage.fir@878.4]
  wire [3:0] _T_542; // @[Lookup.scala 11:37:Sodor3Stage.fir@879.4]
  wire [3:0] _T_543; // @[Lookup.scala 11:37:Sodor3Stage.fir@880.4]
  wire [3:0] _T_544; // @[Lookup.scala 11:37:Sodor3Stage.fir@881.4]
  wire [3:0] _T_545; // @[Lookup.scala 11:37:Sodor3Stage.fir@882.4]
  wire [3:0] _T_546; // @[Lookup.scala 11:37:Sodor3Stage.fir@883.4]
  wire [3:0] _T_547; // @[Lookup.scala 11:37:Sodor3Stage.fir@884.4]
  wire [3:0] _T_548; // @[Lookup.scala 11:37:Sodor3Stage.fir@885.4]
  wire [3:0] _T_549; // @[Lookup.scala 11:37:Sodor3Stage.fir@886.4]
  wire [3:0] _T_550; // @[Lookup.scala 11:37:Sodor3Stage.fir@887.4]
  wire [3:0] _T_551; // @[Lookup.scala 11:37:Sodor3Stage.fir@888.4]
  wire [3:0] _T_552; // @[Lookup.scala 11:37:Sodor3Stage.fir@889.4]
  wire [3:0] _T_553; // @[Lookup.scala 11:37:Sodor3Stage.fir@890.4]
  wire [3:0] _T_554; // @[Lookup.scala 11:37:Sodor3Stage.fir@891.4]
  wire [3:0] _T_555; // @[Lookup.scala 11:37:Sodor3Stage.fir@892.4]
  wire [3:0] _T_556; // @[Lookup.scala 11:37:Sodor3Stage.fir@893.4]
  wire [3:0] _T_557; // @[Lookup.scala 11:37:Sodor3Stage.fir@894.4]
  wire [3:0] _T_558; // @[Lookup.scala 11:37:Sodor3Stage.fir@895.4]
  wire [3:0] _T_559; // @[Lookup.scala 11:37:Sodor3Stage.fir@896.4]
  wire [3:0] _T_560; // @[Lookup.scala 11:37:Sodor3Stage.fir@897.4]
  wire [3:0] _T_561; // @[Lookup.scala 11:37:Sodor3Stage.fir@898.4]
  wire [3:0] _T_562; // @[Lookup.scala 11:37:Sodor3Stage.fir@899.4]
  wire [3:0] _T_563; // @[Lookup.scala 11:37:Sodor3Stage.fir@900.4]
  wire [3:0] _T_564; // @[Lookup.scala 11:37:Sodor3Stage.fir@901.4]
  wire [3:0] _T_565; // @[Lookup.scala 11:37:Sodor3Stage.fir@902.4]
  wire [3:0] _T_566; // @[Lookup.scala 11:37:Sodor3Stage.fir@903.4]
  wire [3:0] _T_567; // @[Lookup.scala 11:37:Sodor3Stage.fir@904.4]
  wire [3:0] _T_568; // @[Lookup.scala 11:37:Sodor3Stage.fir@905.4]
  wire [3:0] _T_569; // @[Lookup.scala 11:37:Sodor3Stage.fir@906.4]
  wire [3:0] _T_570; // @[Lookup.scala 11:37:Sodor3Stage.fir@907.4]
  wire [3:0] _T_571; // @[Lookup.scala 11:37:Sodor3Stage.fir@908.4]
  wire [3:0] _T_572; // @[Lookup.scala 11:37:Sodor3Stage.fir@909.4]
  wire [3:0] _T_573; // @[Lookup.scala 11:37:Sodor3Stage.fir@910.4]
  wire [3:0] _T_574; // @[Lookup.scala 11:37:Sodor3Stage.fir@911.4]
  wire [3:0] _T_575; // @[Lookup.scala 11:37:Sodor3Stage.fir@912.4]
  wire [3:0] _T_576; // @[Lookup.scala 11:37:Sodor3Stage.fir@913.4]
  wire [3:0] _T_577; // @[Lookup.scala 11:37:Sodor3Stage.fir@914.4]
  wire [3:0] _T_578; // @[Lookup.scala 11:37:Sodor3Stage.fir@915.4]
  wire [3:0] _T_579; // @[Lookup.scala 11:37:Sodor3Stage.fir@916.4]
  wire [1:0] _T_587; // @[Lookup.scala 11:37:Sodor3Stage.fir@925.4]
  wire [1:0] _T_588; // @[Lookup.scala 11:37:Sodor3Stage.fir@926.4]
  wire [1:0] _T_589; // @[Lookup.scala 11:37:Sodor3Stage.fir@927.4]
  wire [1:0] _T_590; // @[Lookup.scala 11:37:Sodor3Stage.fir@928.4]
  wire [1:0] _T_591; // @[Lookup.scala 11:37:Sodor3Stage.fir@929.4]
  wire [1:0] _T_592; // @[Lookup.scala 11:37:Sodor3Stage.fir@930.4]
  wire [1:0] _T_593; // @[Lookup.scala 11:37:Sodor3Stage.fir@931.4]
  wire [1:0] _T_594; // @[Lookup.scala 11:37:Sodor3Stage.fir@932.4]
  wire [1:0] _T_595; // @[Lookup.scala 11:37:Sodor3Stage.fir@933.4]
  wire [1:0] _T_596; // @[Lookup.scala 11:37:Sodor3Stage.fir@934.4]
  wire [1:0] _T_597; // @[Lookup.scala 11:37:Sodor3Stage.fir@935.4]
  wire [1:0] _T_598; // @[Lookup.scala 11:37:Sodor3Stage.fir@936.4]
  wire [1:0] _T_599; // @[Lookup.scala 11:37:Sodor3Stage.fir@937.4]
  wire [1:0] _T_600; // @[Lookup.scala 11:37:Sodor3Stage.fir@938.4]
  wire [1:0] _T_601; // @[Lookup.scala 11:37:Sodor3Stage.fir@939.4]
  wire [1:0] _T_602; // @[Lookup.scala 11:37:Sodor3Stage.fir@940.4]
  wire [1:0] _T_603; // @[Lookup.scala 11:37:Sodor3Stage.fir@941.4]
  wire [1:0] _T_604; // @[Lookup.scala 11:37:Sodor3Stage.fir@942.4]
  wire [1:0] _T_605; // @[Lookup.scala 11:37:Sodor3Stage.fir@943.4]
  wire [1:0] _T_606; // @[Lookup.scala 11:37:Sodor3Stage.fir@944.4]
  wire [1:0] _T_607; // @[Lookup.scala 11:37:Sodor3Stage.fir@945.4]
  wire [1:0] _T_608; // @[Lookup.scala 11:37:Sodor3Stage.fir@946.4]
  wire [1:0] _T_609; // @[Lookup.scala 11:37:Sodor3Stage.fir@947.4]
  wire [1:0] _T_610; // @[Lookup.scala 11:37:Sodor3Stage.fir@948.4]
  wire [1:0] _T_611; // @[Lookup.scala 11:37:Sodor3Stage.fir@949.4]
  wire [1:0] _T_612; // @[Lookup.scala 11:37:Sodor3Stage.fir@950.4]
  wire [1:0] _T_613; // @[Lookup.scala 11:37:Sodor3Stage.fir@951.4]
  wire [1:0] _T_614; // @[Lookup.scala 11:37:Sodor3Stage.fir@952.4]
  wire [1:0] _T_615; // @[Lookup.scala 11:37:Sodor3Stage.fir@953.4]
  wire [1:0] _T_616; // @[Lookup.scala 11:37:Sodor3Stage.fir@954.4]
  wire [1:0] _T_617; // @[Lookup.scala 11:37:Sodor3Stage.fir@955.4]
  wire [1:0] _T_618; // @[Lookup.scala 11:37:Sodor3Stage.fir@956.4]
  wire [1:0] _T_619; // @[Lookup.scala 11:37:Sodor3Stage.fir@957.4]
  wire [1:0] _T_620; // @[Lookup.scala 11:37:Sodor3Stage.fir@958.4]
  wire [1:0] _T_621; // @[Lookup.scala 11:37:Sodor3Stage.fir@959.4]
  wire [1:0] _T_622; // @[Lookup.scala 11:37:Sodor3Stage.fir@960.4]
  wire [1:0] _T_623; // @[Lookup.scala 11:37:Sodor3Stage.fir@961.4]
  wire [1:0] _T_624; // @[Lookup.scala 11:37:Sodor3Stage.fir@962.4]
  wire [1:0] _T_625; // @[Lookup.scala 11:37:Sodor3Stage.fir@963.4]
  wire [1:0] _T_626; // @[Lookup.scala 11:37:Sodor3Stage.fir@964.4]
  wire [1:0] _T_627; // @[Lookup.scala 11:37:Sodor3Stage.fir@965.4]
  wire [1:0] _T_628; // @[Lookup.scala 11:37:Sodor3Stage.fir@966.4]
  wire  _T_637; // @[Lookup.scala 11:37:Sodor3Stage.fir@976.4]
  wire  _T_638; // @[Lookup.scala 11:37:Sodor3Stage.fir@977.4]
  wire  _T_639; // @[Lookup.scala 11:37:Sodor3Stage.fir@978.4]
  wire  _T_640; // @[Lookup.scala 11:37:Sodor3Stage.fir@979.4]
  wire  _T_641; // @[Lookup.scala 11:37:Sodor3Stage.fir@980.4]
  wire  _T_642; // @[Lookup.scala 11:37:Sodor3Stage.fir@981.4]
  wire  _T_643; // @[Lookup.scala 11:37:Sodor3Stage.fir@982.4]
  wire  _T_644; // @[Lookup.scala 11:37:Sodor3Stage.fir@983.4]
  wire  _T_645; // @[Lookup.scala 11:37:Sodor3Stage.fir@984.4]
  wire  _T_646; // @[Lookup.scala 11:37:Sodor3Stage.fir@985.4]
  wire  _T_647; // @[Lookup.scala 11:37:Sodor3Stage.fir@986.4]
  wire  _T_648; // @[Lookup.scala 11:37:Sodor3Stage.fir@987.4]
  wire  _T_649; // @[Lookup.scala 11:37:Sodor3Stage.fir@988.4]
  wire  _T_650; // @[Lookup.scala 11:37:Sodor3Stage.fir@989.4]
  wire  _T_651; // @[Lookup.scala 11:37:Sodor3Stage.fir@990.4]
  wire  _T_652; // @[Lookup.scala 11:37:Sodor3Stage.fir@991.4]
  wire  _T_653; // @[Lookup.scala 11:37:Sodor3Stage.fir@992.4]
  wire  _T_654; // @[Lookup.scala 11:37:Sodor3Stage.fir@993.4]
  wire  _T_655; // @[Lookup.scala 11:37:Sodor3Stage.fir@994.4]
  wire  _T_656; // @[Lookup.scala 11:37:Sodor3Stage.fir@995.4]
  wire  _T_657; // @[Lookup.scala 11:37:Sodor3Stage.fir@996.4]
  wire  _T_658; // @[Lookup.scala 11:37:Sodor3Stage.fir@997.4]
  wire  _T_659; // @[Lookup.scala 11:37:Sodor3Stage.fir@998.4]
  wire  _T_660; // @[Lookup.scala 11:37:Sodor3Stage.fir@999.4]
  wire  _T_661; // @[Lookup.scala 11:37:Sodor3Stage.fir@1000.4]
  wire  _T_662; // @[Lookup.scala 11:37:Sodor3Stage.fir@1001.4]
  wire  _T_663; // @[Lookup.scala 11:37:Sodor3Stage.fir@1002.4]
  wire  _T_664; // @[Lookup.scala 11:37:Sodor3Stage.fir@1003.4]
  wire  _T_665; // @[Lookup.scala 11:37:Sodor3Stage.fir@1004.4]
  wire  _T_666; // @[Lookup.scala 11:37:Sodor3Stage.fir@1005.4]
  wire  _T_667; // @[Lookup.scala 11:37:Sodor3Stage.fir@1006.4]
  wire  _T_668; // @[Lookup.scala 11:37:Sodor3Stage.fir@1007.4]
  wire  _T_669; // @[Lookup.scala 11:37:Sodor3Stage.fir@1008.4]
  wire  _T_670; // @[Lookup.scala 11:37:Sodor3Stage.fir@1009.4]
  wire  _T_671; // @[Lookup.scala 11:37:Sodor3Stage.fir@1010.4]
  wire  _T_672; // @[Lookup.scala 11:37:Sodor3Stage.fir@1011.4]
  wire  _T_673; // @[Lookup.scala 11:37:Sodor3Stage.fir@1012.4]
  wire  _T_674; // @[Lookup.scala 11:37:Sodor3Stage.fir@1013.4]
  wire  _T_675; // @[Lookup.scala 11:37:Sodor3Stage.fir@1014.4]
  wire  _T_676; // @[Lookup.scala 11:37:Sodor3Stage.fir@1015.4]
  wire  _T_677; // @[Lookup.scala 11:37:Sodor3Stage.fir@1016.4]
  wire  cs0_2; // @[Lookup.scala 11:37:Sodor3Stage.fir@1017.4]
  wire  _T_699; // @[Lookup.scala 11:37:Sodor3Stage.fir@1039.4]
  wire  _T_700; // @[Lookup.scala 11:37:Sodor3Stage.fir@1040.4]
  wire  _T_701; // @[Lookup.scala 11:37:Sodor3Stage.fir@1041.4]
  wire  _T_702; // @[Lookup.scala 11:37:Sodor3Stage.fir@1042.4]
  wire  _T_703; // @[Lookup.scala 11:37:Sodor3Stage.fir@1043.4]
  wire  _T_704; // @[Lookup.scala 11:37:Sodor3Stage.fir@1044.4]
  wire  _T_705; // @[Lookup.scala 11:37:Sodor3Stage.fir@1045.4]
  wire  _T_706; // @[Lookup.scala 11:37:Sodor3Stage.fir@1046.4]
  wire  _T_707; // @[Lookup.scala 11:37:Sodor3Stage.fir@1047.4]
  wire  _T_708; // @[Lookup.scala 11:37:Sodor3Stage.fir@1048.4]
  wire  _T_709; // @[Lookup.scala 11:37:Sodor3Stage.fir@1049.4]
  wire  _T_710; // @[Lookup.scala 11:37:Sodor3Stage.fir@1050.4]
  wire  _T_711; // @[Lookup.scala 11:37:Sodor3Stage.fir@1051.4]
  wire  _T_712; // @[Lookup.scala 11:37:Sodor3Stage.fir@1052.4]
  wire  _T_713; // @[Lookup.scala 11:37:Sodor3Stage.fir@1053.4]
  wire  _T_714; // @[Lookup.scala 11:37:Sodor3Stage.fir@1054.4]
  wire  _T_715; // @[Lookup.scala 11:37:Sodor3Stage.fir@1055.4]
  wire  _T_716; // @[Lookup.scala 11:37:Sodor3Stage.fir@1056.4]
  wire  _T_717; // @[Lookup.scala 11:37:Sodor3Stage.fir@1057.4]
  wire  _T_718; // @[Lookup.scala 11:37:Sodor3Stage.fir@1058.4]
  wire  _T_719; // @[Lookup.scala 11:37:Sodor3Stage.fir@1059.4]
  wire  _T_720; // @[Lookup.scala 11:37:Sodor3Stage.fir@1060.4]
  wire  _T_721; // @[Lookup.scala 11:37:Sodor3Stage.fir@1061.4]
  wire  _T_722; // @[Lookup.scala 11:37:Sodor3Stage.fir@1062.4]
  wire  _T_723; // @[Lookup.scala 11:37:Sodor3Stage.fir@1063.4]
  wire  _T_724; // @[Lookup.scala 11:37:Sodor3Stage.fir@1064.4]
  wire  _T_725; // @[Lookup.scala 11:37:Sodor3Stage.fir@1065.4]
  wire  _T_726; // @[Lookup.scala 11:37:Sodor3Stage.fir@1066.4]
  wire  _T_819; // @[Lookup.scala 11:37:Sodor3Stage.fir@1161.4]
  wire  _T_820; // @[Lookup.scala 11:37:Sodor3Stage.fir@1162.4]
  wire  _T_821; // @[Lookup.scala 11:37:Sodor3Stage.fir@1163.4]
  wire  _T_822; // @[Lookup.scala 11:37:Sodor3Stage.fir@1164.4]
  wire  _T_823; // @[Lookup.scala 11:37:Sodor3Stage.fir@1165.4]
  wire  _T_824; // @[Lookup.scala 11:37:Sodor3Stage.fir@1166.4]
  wire [2:0] _T_867; // @[Lookup.scala 11:37:Sodor3Stage.fir@1210.4]
  wire [2:0] _T_868; // @[Lookup.scala 11:37:Sodor3Stage.fir@1211.4]
  wire [2:0] _T_869; // @[Lookup.scala 11:37:Sodor3Stage.fir@1212.4]
  wire [2:0] _T_870; // @[Lookup.scala 11:37:Sodor3Stage.fir@1213.4]
  wire [2:0] _T_871; // @[Lookup.scala 11:37:Sodor3Stage.fir@1214.4]
  wire [2:0] _T_872; // @[Lookup.scala 11:37:Sodor3Stage.fir@1215.4]
  wire [2:0] _T_873; // @[Lookup.scala 11:37:Sodor3Stage.fir@1216.4]
  wire [2:0] _T_876; // @[Lookup.scala 11:37:Sodor3Stage.fir@1220.4]
  wire [2:0] _T_877; // @[Lookup.scala 11:37:Sodor3Stage.fir@1221.4]
  wire [2:0] _T_878; // @[Lookup.scala 11:37:Sodor3Stage.fir@1222.4]
  wire [2:0] _T_879; // @[Lookup.scala 11:37:Sodor3Stage.fir@1223.4]
  wire [2:0] _T_880; // @[Lookup.scala 11:37:Sodor3Stage.fir@1224.4]
  wire [2:0] _T_881; // @[Lookup.scala 11:37:Sodor3Stage.fir@1225.4]
  wire [2:0] _T_882; // @[Lookup.scala 11:37:Sodor3Stage.fir@1226.4]
  wire [2:0] _T_883; // @[Lookup.scala 11:37:Sodor3Stage.fir@1227.4]
  wire [2:0] _T_884; // @[Lookup.scala 11:37:Sodor3Stage.fir@1228.4]
  wire [2:0] _T_885; // @[Lookup.scala 11:37:Sodor3Stage.fir@1229.4]
  wire [2:0] _T_886; // @[Lookup.scala 11:37:Sodor3Stage.fir@1230.4]
  wire [2:0] _T_887; // @[Lookup.scala 11:37:Sodor3Stage.fir@1231.4]
  wire [2:0] _T_888; // @[Lookup.scala 11:37:Sodor3Stage.fir@1232.4]
  wire [2:0] _T_889; // @[Lookup.scala 11:37:Sodor3Stage.fir@1233.4]
  wire [2:0] _T_890; // @[Lookup.scala 11:37:Sodor3Stage.fir@1234.4]
  wire [2:0] _T_891; // @[Lookup.scala 11:37:Sodor3Stage.fir@1235.4]
  wire [2:0] _T_892; // @[Lookup.scala 11:37:Sodor3Stage.fir@1236.4]
  wire [2:0] _T_893; // @[Lookup.scala 11:37:Sodor3Stage.fir@1237.4]
  wire [2:0] _T_894; // @[Lookup.scala 11:37:Sodor3Stage.fir@1238.4]
  wire [2:0] _T_895; // @[Lookup.scala 11:37:Sodor3Stage.fir@1239.4]
  wire [2:0] _T_896; // @[Lookup.scala 11:37:Sodor3Stage.fir@1240.4]
  wire [2:0] _T_897; // @[Lookup.scala 11:37:Sodor3Stage.fir@1241.4]
  wire [2:0] _T_898; // @[Lookup.scala 11:37:Sodor3Stage.fir@1242.4]
  wire [2:0] _T_899; // @[Lookup.scala 11:37:Sodor3Stage.fir@1243.4]
  wire [2:0] _T_900; // @[Lookup.scala 11:37:Sodor3Stage.fir@1244.4]
  wire [2:0] _T_901; // @[Lookup.scala 11:37:Sodor3Stage.fir@1245.4]
  wire [2:0] _T_902; // @[Lookup.scala 11:37:Sodor3Stage.fir@1246.4]
  wire [2:0] _T_903; // @[Lookup.scala 11:37:Sodor3Stage.fir@1247.4]
  wire [2:0] _T_904; // @[Lookup.scala 11:37:Sodor3Stage.fir@1248.4]
  wire [2:0] _T_905; // @[Lookup.scala 11:37:Sodor3Stage.fir@1249.4]
  wire [2:0] _T_906; // @[Lookup.scala 11:37:Sodor3Stage.fir@1250.4]
  wire [2:0] _T_907; // @[Lookup.scala 11:37:Sodor3Stage.fir@1251.4]
  wire [2:0] _T_908; // @[Lookup.scala 11:37:Sodor3Stage.fir@1252.4]
  wire [2:0] _T_909; // @[Lookup.scala 11:37:Sodor3Stage.fir@1253.4]
  wire [2:0] _T_910; // @[Lookup.scala 11:37:Sodor3Stage.fir@1254.4]
  wire [2:0] _T_911; // @[Lookup.scala 11:37:Sodor3Stage.fir@1255.4]
  wire [2:0] _T_912; // @[Lookup.scala 11:37:Sodor3Stage.fir@1256.4]
  wire [2:0] _T_913; // @[Lookup.scala 11:37:Sodor3Stage.fir@1257.4]
  wire [2:0] _T_914; // @[Lookup.scala 11:37:Sodor3Stage.fir@1258.4]
  wire [2:0] _T_915; // @[Lookup.scala 11:37:Sodor3Stage.fir@1259.4]
  wire [2:0] _T_916; // @[Lookup.scala 11:37:Sodor3Stage.fir@1260.4]
  wire [2:0] _T_917; // @[Lookup.scala 11:37:Sodor3Stage.fir@1261.4]
  wire [2:0] _T_918; // @[Lookup.scala 11:37:Sodor3Stage.fir@1262.4]
  wire [2:0] _T_919; // @[Lookup.scala 11:37:Sodor3Stage.fir@1263.4]
  wire [2:0] _T_920; // @[Lookup.scala 11:37:Sodor3Stage.fir@1264.4]
  wire [2:0] _T_921; // @[Lookup.scala 11:37:Sodor3Stage.fir@1265.4]
  wire [2:0] _T_922; // @[Lookup.scala 11:37:Sodor3Stage.fir@1266.4]
  wire [2:0] cs0_7; // @[Lookup.scala 11:37:Sodor3Stage.fir@1267.4]
  wire  _T_973; // @[cpath.scala 138:37:Sodor3Stage.fir@1319.4]
  wire  _T_974; // @[cpath.scala 139:37:Sodor3Stage.fir@1320.4]
  wire  _T_976; // @[cpath.scala 139:54:Sodor3Stage.fir@1321.4]
  wire [2:0] _T_977; // @[cpath.scala 139:53:Sodor3Stage.fir@1322.4]
  wire  _T_978; // @[cpath.scala 140:37:Sodor3Stage.fir@1323.4]
  wire [2:0] _T_979; // @[cpath.scala 140:53:Sodor3Stage.fir@1324.4]
  wire  _T_980; // @[cpath.scala 141:37:Sodor3Stage.fir@1325.4]
  wire  _T_982; // @[cpath.scala 141:54:Sodor3Stage.fir@1326.4]
  wire [2:0] _T_983; // @[cpath.scala 141:53:Sodor3Stage.fir@1327.4]
  wire  _T_984; // @[cpath.scala 142:37:Sodor3Stage.fir@1328.4]
  wire  _T_986; // @[cpath.scala 142:54:Sodor3Stage.fir@1329.4]
  wire [2:0] _T_987; // @[cpath.scala 142:53:Sodor3Stage.fir@1330.4]
  wire  _T_988; // @[cpath.scala 143:37:Sodor3Stage.fir@1331.4]
  wire [2:0] _T_989; // @[cpath.scala 143:53:Sodor3Stage.fir@1332.4]
  wire  _T_990; // @[cpath.scala 144:37:Sodor3Stage.fir@1333.4]
  wire [2:0] _T_991; // @[cpath.scala 144:53:Sodor3Stage.fir@1334.4]
  wire  _T_992; // @[cpath.scala 145:37:Sodor3Stage.fir@1335.4]
  wire  _T_993; // @[cpath.scala 146:37:Sodor3Stage.fir@1336.4]
  wire [2:0] _T_994; // @[cpath.scala 146:25:Sodor3Stage.fir@1337.4]
  wire [2:0] _T_995; // @[cpath.scala 145:25:Sodor3Stage.fir@1338.4]
  wire [2:0] _T_996; // @[cpath.scala 144:25:Sodor3Stage.fir@1339.4]
  wire [2:0] _T_997; // @[cpath.scala 143:25:Sodor3Stage.fir@1340.4]
  wire [2:0] _T_998; // @[cpath.scala 142:25:Sodor3Stage.fir@1341.4]
  wire [2:0] _T_999; // @[cpath.scala 141:25:Sodor3Stage.fir@1342.4]
  wire [2:0] _T_1000; // @[cpath.scala 140:25:Sodor3Stage.fir@1343.4]
  wire [2:0] _T_1001; // @[cpath.scala 139:25:Sodor3Stage.fir@1344.4]
  wire [2:0] _T_1002; // @[cpath.scala 138:25:Sodor3Stage.fir@1345.4]
  wire  take_evec; // @[cpath.scala 179:51:Sodor3Stage.fir@1385.4]
  wire [2:0] ctrl_pc_sel; // @[cpath.scala 137:25:Sodor3Stage.fir@1346.4]
  wire  _T_1003; // @[cpath.scala 150:39:Sodor3Stage.fir@1347.4]
  wire  _T_1005; // @[cpath.scala 150:25:Sodor3Stage.fir@1348.4]
  wire  _T_1009; // @[cpath.scala 159:29:Sodor3Stage.fir@1359.4]
  wire [4:0] rs1_addr; // @[cpath.scala 162:41:Sodor3Stage.fir@1365.4]
  wire  _T_1014; // @[cpath.scala 163:30:Sodor3Stage.fir@1366.4]
  wire  _T_1015; // @[cpath.scala 163:54:Sodor3Stage.fir@1367.4]
  wire  _T_1016; // @[cpath.scala 163:40:Sodor3Stage.fir@1368.4]
  wire  _T_1018; // @[cpath.scala 163:77:Sodor3Stage.fir@1369.4]
  wire  csr_ren; // @[cpath.scala 163:65:Sodor3Stage.fir@1370.4]
  wire [2:0] csr_cmd; // @[cpath.scala 164:21:Sodor3Stage.fir@1371.4]
  wire  _T_1025; // @[cpath.scala 178:24:Sodor3Stage.fir@1380.4]
  assign _T_88 = io_imem_resp_bits_inst & 32'h707f; // @[Lookup.scala 9:38:Sodor3Stage.fir@518.4]
  assign _T_89 = 32'h2003 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@519.4]
  assign _T_93 = 32'h3 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@521.4]
  assign _T_97 = 32'h4003 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@523.4]
  assign _T_101 = 32'h1003 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@525.4]
  assign _T_105 = 32'h5003 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@527.4]
  assign _T_109 = 32'h2023 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@529.4]
  assign _T_113 = 32'h23 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@531.4]
  assign _T_117 = 32'h1023 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@533.4]
  assign _T_120 = io_imem_resp_bits_inst & 32'h7f; // @[Lookup.scala 9:38:Sodor3Stage.fir@534.4]
  assign _T_121 = 32'h17 == _T_120; // @[Lookup.scala 9:38:Sodor3Stage.fir@535.4]
  assign _T_125 = 32'h37 == _T_120; // @[Lookup.scala 9:38:Sodor3Stage.fir@537.4]
  assign _T_129 = 32'h13 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@539.4]
  assign _T_133 = 32'h7013 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@541.4]
  assign _T_137 = 32'h6013 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@543.4]
  assign _T_141 = 32'h4013 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@545.4]
  assign _T_145 = 32'h2013 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@547.4]
  assign _T_149 = 32'h3013 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@549.4]
  assign _T_152 = io_imem_resp_bits_inst & 32'hfc00707f; // @[Lookup.scala 9:38:Sodor3Stage.fir@550.4]
  assign _T_153 = 32'h1013 == _T_152; // @[Lookup.scala 9:38:Sodor3Stage.fir@551.4]
  assign _T_157 = 32'h40005013 == _T_152; // @[Lookup.scala 9:38:Sodor3Stage.fir@553.4]
  assign _T_161 = 32'h5013 == _T_152; // @[Lookup.scala 9:38:Sodor3Stage.fir@555.4]
  assign _T_164 = io_imem_resp_bits_inst & 32'hfe00707f; // @[Lookup.scala 9:38:Sodor3Stage.fir@556.4]
  assign _T_165 = 32'h1033 == _T_164; // @[Lookup.scala 9:38:Sodor3Stage.fir@557.4]
  assign _T_169 = 32'h33 == _T_164; // @[Lookup.scala 9:38:Sodor3Stage.fir@559.4]
  assign _T_173 = 32'h40000033 == _T_164; // @[Lookup.scala 9:38:Sodor3Stage.fir@561.4]
  assign _T_177 = 32'h2033 == _T_164; // @[Lookup.scala 9:38:Sodor3Stage.fir@563.4]
  assign _T_181 = 32'h3033 == _T_164; // @[Lookup.scala 9:38:Sodor3Stage.fir@565.4]
  assign _T_185 = 32'h7033 == _T_164; // @[Lookup.scala 9:38:Sodor3Stage.fir@567.4]
  assign _T_189 = 32'h6033 == _T_164; // @[Lookup.scala 9:38:Sodor3Stage.fir@569.4]
  assign _T_193 = 32'h4033 == _T_164; // @[Lookup.scala 9:38:Sodor3Stage.fir@571.4]
  assign _T_197 = 32'h40005033 == _T_164; // @[Lookup.scala 9:38:Sodor3Stage.fir@573.4]
  assign _T_201 = 32'h5033 == _T_164; // @[Lookup.scala 9:38:Sodor3Stage.fir@575.4]
  assign _T_205 = 32'h6f == _T_120; // @[Lookup.scala 9:38:Sodor3Stage.fir@577.4]
  assign _T_209 = 32'h67 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@579.4]
  assign _T_213 = 32'h63 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@581.4]
  assign _T_217 = 32'h1063 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@583.4]
  assign _T_221 = 32'h5063 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@585.4]
  assign _T_225 = 32'h7063 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@587.4]
  assign _T_229 = 32'h4063 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@589.4]
  assign _T_233 = 32'h6063 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@591.4]
  assign _T_237 = 32'h5073 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@593.4]
  assign _T_241 = 32'h6073 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@595.4]
  assign _T_245 = 32'h1073 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@597.4]
  assign _T_249 = 32'h2073 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@599.4]
  assign _T_253 = 32'h3073 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@601.4]
  assign _T_257 = 32'h7073 == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@603.4]
  assign _T_261 = 32'h73 == io_imem_resp_bits_inst; // @[Lookup.scala 9:38:Sodor3Stage.fir@605.4]
  assign _T_265 = 32'h30200073 == io_imem_resp_bits_inst; // @[Lookup.scala 9:38:Sodor3Stage.fir@607.4]
  assign _T_269 = 32'h7b200073 == io_imem_resp_bits_inst; // @[Lookup.scala 9:38:Sodor3Stage.fir@609.4]
  assign _T_273 = 32'h100073 == io_imem_resp_bits_inst; // @[Lookup.scala 9:38:Sodor3Stage.fir@611.4]
  assign _T_277 = 32'h10500073 == io_imem_resp_bits_inst; // @[Lookup.scala 9:38:Sodor3Stage.fir@613.4]
  assign _T_281 = 32'h100f == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@615.4]
  assign _T_285 = 32'hf == _T_88; // @[Lookup.scala 9:38:Sodor3Stage.fir@617.4]
  assign _T_287 = _T_281 ? 1'h1 : _T_285; // @[Lookup.scala 11:37:Sodor3Stage.fir@619.4]
  assign _T_288 = _T_277 ? 1'h1 : _T_287; // @[Lookup.scala 11:37:Sodor3Stage.fir@620.4]
  assign _T_289 = _T_273 ? 1'h1 : _T_288; // @[Lookup.scala 11:37:Sodor3Stage.fir@621.4]
  assign _T_290 = _T_269 ? 1'h1 : _T_289; // @[Lookup.scala 11:37:Sodor3Stage.fir@622.4]
  assign _T_291 = _T_265 ? 1'h1 : _T_290; // @[Lookup.scala 11:37:Sodor3Stage.fir@623.4]
  assign _T_292 = _T_261 ? 1'h1 : _T_291; // @[Lookup.scala 11:37:Sodor3Stage.fir@624.4]
  assign _T_293 = _T_257 ? 1'h1 : _T_292; // @[Lookup.scala 11:37:Sodor3Stage.fir@625.4]
  assign _T_294 = _T_253 ? 1'h1 : _T_293; // @[Lookup.scala 11:37:Sodor3Stage.fir@626.4]
  assign _T_295 = _T_249 ? 1'h1 : _T_294; // @[Lookup.scala 11:37:Sodor3Stage.fir@627.4]
  assign _T_296 = _T_245 ? 1'h1 : _T_295; // @[Lookup.scala 11:37:Sodor3Stage.fir@628.4]
  assign _T_297 = _T_241 ? 1'h1 : _T_296; // @[Lookup.scala 11:37:Sodor3Stage.fir@629.4]
  assign _T_298 = _T_237 ? 1'h1 : _T_297; // @[Lookup.scala 11:37:Sodor3Stage.fir@630.4]
  assign _T_299 = _T_233 ? 1'h1 : _T_298; // @[Lookup.scala 11:37:Sodor3Stage.fir@631.4]
  assign _T_300 = _T_229 ? 1'h1 : _T_299; // @[Lookup.scala 11:37:Sodor3Stage.fir@632.4]
  assign _T_301 = _T_225 ? 1'h1 : _T_300; // @[Lookup.scala 11:37:Sodor3Stage.fir@633.4]
  assign _T_302 = _T_221 ? 1'h1 : _T_301; // @[Lookup.scala 11:37:Sodor3Stage.fir@634.4]
  assign _T_303 = _T_217 ? 1'h1 : _T_302; // @[Lookup.scala 11:37:Sodor3Stage.fir@635.4]
  assign _T_304 = _T_213 ? 1'h1 : _T_303; // @[Lookup.scala 11:37:Sodor3Stage.fir@636.4]
  assign _T_305 = _T_209 ? 1'h1 : _T_304; // @[Lookup.scala 11:37:Sodor3Stage.fir@637.4]
  assign _T_306 = _T_205 ? 1'h1 : _T_305; // @[Lookup.scala 11:37:Sodor3Stage.fir@638.4]
  assign _T_307 = _T_201 ? 1'h1 : _T_306; // @[Lookup.scala 11:37:Sodor3Stage.fir@639.4]
  assign _T_308 = _T_197 ? 1'h1 : _T_307; // @[Lookup.scala 11:37:Sodor3Stage.fir@640.4]
  assign _T_309 = _T_193 ? 1'h1 : _T_308; // @[Lookup.scala 11:37:Sodor3Stage.fir@641.4]
  assign _T_310 = _T_189 ? 1'h1 : _T_309; // @[Lookup.scala 11:37:Sodor3Stage.fir@642.4]
  assign _T_311 = _T_185 ? 1'h1 : _T_310; // @[Lookup.scala 11:37:Sodor3Stage.fir@643.4]
  assign _T_312 = _T_181 ? 1'h1 : _T_311; // @[Lookup.scala 11:37:Sodor3Stage.fir@644.4]
  assign _T_313 = _T_177 ? 1'h1 : _T_312; // @[Lookup.scala 11:37:Sodor3Stage.fir@645.4]
  assign _T_314 = _T_173 ? 1'h1 : _T_313; // @[Lookup.scala 11:37:Sodor3Stage.fir@646.4]
  assign _T_315 = _T_169 ? 1'h1 : _T_314; // @[Lookup.scala 11:37:Sodor3Stage.fir@647.4]
  assign _T_316 = _T_165 ? 1'h1 : _T_315; // @[Lookup.scala 11:37:Sodor3Stage.fir@648.4]
  assign _T_317 = _T_161 ? 1'h1 : _T_316; // @[Lookup.scala 11:37:Sodor3Stage.fir@649.4]
  assign _T_318 = _T_157 ? 1'h1 : _T_317; // @[Lookup.scala 11:37:Sodor3Stage.fir@650.4]
  assign _T_319 = _T_153 ? 1'h1 : _T_318; // @[Lookup.scala 11:37:Sodor3Stage.fir@651.4]
  assign _T_320 = _T_149 ? 1'h1 : _T_319; // @[Lookup.scala 11:37:Sodor3Stage.fir@652.4]
  assign _T_321 = _T_145 ? 1'h1 : _T_320; // @[Lookup.scala 11:37:Sodor3Stage.fir@653.4]
  assign _T_322 = _T_141 ? 1'h1 : _T_321; // @[Lookup.scala 11:37:Sodor3Stage.fir@654.4]
  assign _T_323 = _T_137 ? 1'h1 : _T_322; // @[Lookup.scala 11:37:Sodor3Stage.fir@655.4]
  assign _T_324 = _T_133 ? 1'h1 : _T_323; // @[Lookup.scala 11:37:Sodor3Stage.fir@656.4]
  assign _T_325 = _T_129 ? 1'h1 : _T_324; // @[Lookup.scala 11:37:Sodor3Stage.fir@657.4]
  assign _T_326 = _T_125 ? 1'h1 : _T_325; // @[Lookup.scala 11:37:Sodor3Stage.fir@658.4]
  assign _T_327 = _T_121 ? 1'h1 : _T_326; // @[Lookup.scala 11:37:Sodor3Stage.fir@659.4]
  assign _T_328 = _T_117 ? 1'h1 : _T_327; // @[Lookup.scala 11:37:Sodor3Stage.fir@660.4]
  assign _T_329 = _T_113 ? 1'h1 : _T_328; // @[Lookup.scala 11:37:Sodor3Stage.fir@661.4]
  assign _T_330 = _T_109 ? 1'h1 : _T_329; // @[Lookup.scala 11:37:Sodor3Stage.fir@662.4]
  assign _T_331 = _T_105 ? 1'h1 : _T_330; // @[Lookup.scala 11:37:Sodor3Stage.fir@663.4]
  assign _T_332 = _T_101 ? 1'h1 : _T_331; // @[Lookup.scala 11:37:Sodor3Stage.fir@664.4]
  assign _T_333 = _T_97 ? 1'h1 : _T_332; // @[Lookup.scala 11:37:Sodor3Stage.fir@665.4]
  assign _T_334 = _T_93 ? 1'h1 : _T_333; // @[Lookup.scala 11:37:Sodor3Stage.fir@666.4]
  assign cs_inst_val = _T_89 ? 1'h1 : _T_334; // @[Lookup.scala 11:37:Sodor3Stage.fir@667.4]
  assign _T_348 = _T_233 ? 4'h6 : 4'h0; // @[Lookup.scala 11:37:Sodor3Stage.fir@681.4]
  assign _T_349 = _T_229 ? 4'h5 : _T_348; // @[Lookup.scala 11:37:Sodor3Stage.fir@682.4]
  assign _T_350 = _T_225 ? 4'h4 : _T_349; // @[Lookup.scala 11:37:Sodor3Stage.fir@683.4]
  assign _T_351 = _T_221 ? 4'h3 : _T_350; // @[Lookup.scala 11:37:Sodor3Stage.fir@684.4]
  assign _T_352 = _T_217 ? 4'h1 : _T_351; // @[Lookup.scala 11:37:Sodor3Stage.fir@685.4]
  assign _T_353 = _T_213 ? 4'h2 : _T_352; // @[Lookup.scala 11:37:Sodor3Stage.fir@686.4]
  assign _T_354 = _T_209 ? 4'h8 : _T_353; // @[Lookup.scala 11:37:Sodor3Stage.fir@687.4]
  assign _T_355 = _T_205 ? 4'h7 : _T_354; // @[Lookup.scala 11:37:Sodor3Stage.fir@688.4]
  assign _T_356 = _T_201 ? 4'h0 : _T_355; // @[Lookup.scala 11:37:Sodor3Stage.fir@689.4]
  assign _T_357 = _T_197 ? 4'h0 : _T_356; // @[Lookup.scala 11:37:Sodor3Stage.fir@690.4]
  assign _T_358 = _T_193 ? 4'h0 : _T_357; // @[Lookup.scala 11:37:Sodor3Stage.fir@691.4]
  assign _T_359 = _T_189 ? 4'h0 : _T_358; // @[Lookup.scala 11:37:Sodor3Stage.fir@692.4]
  assign _T_360 = _T_185 ? 4'h0 : _T_359; // @[Lookup.scala 11:37:Sodor3Stage.fir@693.4]
  assign _T_361 = _T_181 ? 4'h0 : _T_360; // @[Lookup.scala 11:37:Sodor3Stage.fir@694.4]
  assign _T_362 = _T_177 ? 4'h0 : _T_361; // @[Lookup.scala 11:37:Sodor3Stage.fir@695.4]
  assign _T_363 = _T_173 ? 4'h0 : _T_362; // @[Lookup.scala 11:37:Sodor3Stage.fir@696.4]
  assign _T_364 = _T_169 ? 4'h0 : _T_363; // @[Lookup.scala 11:37:Sodor3Stage.fir@697.4]
  assign _T_365 = _T_165 ? 4'h0 : _T_364; // @[Lookup.scala 11:37:Sodor3Stage.fir@698.4]
  assign _T_366 = _T_161 ? 4'h0 : _T_365; // @[Lookup.scala 11:37:Sodor3Stage.fir@699.4]
  assign _T_367 = _T_157 ? 4'h0 : _T_366; // @[Lookup.scala 11:37:Sodor3Stage.fir@700.4]
  assign _T_368 = _T_153 ? 4'h0 : _T_367; // @[Lookup.scala 11:37:Sodor3Stage.fir@701.4]
  assign _T_369 = _T_149 ? 4'h0 : _T_368; // @[Lookup.scala 11:37:Sodor3Stage.fir@702.4]
  assign _T_370 = _T_145 ? 4'h0 : _T_369; // @[Lookup.scala 11:37:Sodor3Stage.fir@703.4]
  assign _T_371 = _T_141 ? 4'h0 : _T_370; // @[Lookup.scala 11:37:Sodor3Stage.fir@704.4]
  assign _T_372 = _T_137 ? 4'h0 : _T_371; // @[Lookup.scala 11:37:Sodor3Stage.fir@705.4]
  assign _T_373 = _T_133 ? 4'h0 : _T_372; // @[Lookup.scala 11:37:Sodor3Stage.fir@706.4]
  assign _T_374 = _T_129 ? 4'h0 : _T_373; // @[Lookup.scala 11:37:Sodor3Stage.fir@707.4]
  assign _T_375 = _T_125 ? 4'h0 : _T_374; // @[Lookup.scala 11:37:Sodor3Stage.fir@708.4]
  assign _T_376 = _T_121 ? 4'h0 : _T_375; // @[Lookup.scala 11:37:Sodor3Stage.fir@709.4]
  assign _T_377 = _T_117 ? 4'h0 : _T_376; // @[Lookup.scala 11:37:Sodor3Stage.fir@710.4]
  assign _T_378 = _T_113 ? 4'h0 : _T_377; // @[Lookup.scala 11:37:Sodor3Stage.fir@711.4]
  assign _T_379 = _T_109 ? 4'h0 : _T_378; // @[Lookup.scala 11:37:Sodor3Stage.fir@712.4]
  assign _T_380 = _T_105 ? 4'h0 : _T_379; // @[Lookup.scala 11:37:Sodor3Stage.fir@713.4]
  assign _T_381 = _T_101 ? 4'h0 : _T_380; // @[Lookup.scala 11:37:Sodor3Stage.fir@714.4]
  assign _T_382 = _T_97 ? 4'h0 : _T_381; // @[Lookup.scala 11:37:Sodor3Stage.fir@715.4]
  assign _T_383 = _T_93 ? 4'h0 : _T_382; // @[Lookup.scala 11:37:Sodor3Stage.fir@716.4]
  assign cs_br_type = _T_89 ? 4'h0 : _T_383; // @[Lookup.scala 11:37:Sodor3Stage.fir@717.4]
  assign _T_404 = _T_205 ? 1'h1 : _T_209; // @[Lookup.scala 11:37:Sodor3Stage.fir@738.4]
  assign _T_405 = _T_201 ? 1'h0 : _T_404; // @[Lookup.scala 11:37:Sodor3Stage.fir@739.4]
  assign _T_406 = _T_197 ? 1'h0 : _T_405; // @[Lookup.scala 11:37:Sodor3Stage.fir@740.4]
  assign _T_407 = _T_193 ? 1'h0 : _T_406; // @[Lookup.scala 11:37:Sodor3Stage.fir@741.4]
  assign _T_408 = _T_189 ? 1'h0 : _T_407; // @[Lookup.scala 11:37:Sodor3Stage.fir@742.4]
  assign _T_409 = _T_185 ? 1'h0 : _T_408; // @[Lookup.scala 11:37:Sodor3Stage.fir@743.4]
  assign _T_410 = _T_181 ? 1'h0 : _T_409; // @[Lookup.scala 11:37:Sodor3Stage.fir@744.4]
  assign _T_411 = _T_177 ? 1'h0 : _T_410; // @[Lookup.scala 11:37:Sodor3Stage.fir@745.4]
  assign _T_412 = _T_173 ? 1'h0 : _T_411; // @[Lookup.scala 11:37:Sodor3Stage.fir@746.4]
  assign _T_413 = _T_169 ? 1'h0 : _T_412; // @[Lookup.scala 11:37:Sodor3Stage.fir@747.4]
  assign _T_414 = _T_165 ? 1'h0 : _T_413; // @[Lookup.scala 11:37:Sodor3Stage.fir@748.4]
  assign _T_415 = _T_161 ? 1'h0 : _T_414; // @[Lookup.scala 11:37:Sodor3Stage.fir@749.4]
  assign _T_416 = _T_157 ? 1'h0 : _T_415; // @[Lookup.scala 11:37:Sodor3Stage.fir@750.4]
  assign _T_417 = _T_153 ? 1'h0 : _T_416; // @[Lookup.scala 11:37:Sodor3Stage.fir@751.4]
  assign _T_418 = _T_149 ? 1'h0 : _T_417; // @[Lookup.scala 11:37:Sodor3Stage.fir@752.4]
  assign _T_419 = _T_145 ? 1'h0 : _T_418; // @[Lookup.scala 11:37:Sodor3Stage.fir@753.4]
  assign _T_420 = _T_141 ? 1'h0 : _T_419; // @[Lookup.scala 11:37:Sodor3Stage.fir@754.4]
  assign _T_421 = _T_137 ? 1'h0 : _T_420; // @[Lookup.scala 11:37:Sodor3Stage.fir@755.4]
  assign _T_422 = _T_133 ? 1'h0 : _T_421; // @[Lookup.scala 11:37:Sodor3Stage.fir@756.4]
  assign _T_423 = _T_129 ? 1'h0 : _T_422; // @[Lookup.scala 11:37:Sodor3Stage.fir@757.4]
  assign _T_424 = _T_125 ? 1'h0 : _T_423; // @[Lookup.scala 11:37:Sodor3Stage.fir@758.4]
  assign _T_425 = _T_121 ? 1'h0 : _T_424; // @[Lookup.scala 11:37:Sodor3Stage.fir@759.4]
  assign _T_426 = _T_117 ? 1'h0 : _T_425; // @[Lookup.scala 11:37:Sodor3Stage.fir@760.4]
  assign _T_427 = _T_113 ? 1'h0 : _T_426; // @[Lookup.scala 11:37:Sodor3Stage.fir@761.4]
  assign _T_428 = _T_109 ? 1'h0 : _T_427; // @[Lookup.scala 11:37:Sodor3Stage.fir@762.4]
  assign _T_429 = _T_105 ? 1'h0 : _T_428; // @[Lookup.scala 11:37:Sodor3Stage.fir@763.4]
  assign _T_430 = _T_101 ? 1'h0 : _T_429; // @[Lookup.scala 11:37:Sodor3Stage.fir@764.4]
  assign _T_431 = _T_97 ? 1'h0 : _T_430; // @[Lookup.scala 11:37:Sodor3Stage.fir@765.4]
  assign _T_432 = _T_93 ? 1'h0 : _T_431; // @[Lookup.scala 11:37:Sodor3Stage.fir@766.4]
  assign _T_440 = _T_257 ? 2'h2 : 2'h0; // @[Lookup.scala 11:37:Sodor3Stage.fir@775.4]
  assign _T_441 = _T_253 ? 2'h0 : _T_440; // @[Lookup.scala 11:37:Sodor3Stage.fir@776.4]
  assign _T_442 = _T_249 ? 2'h0 : _T_441; // @[Lookup.scala 11:37:Sodor3Stage.fir@777.4]
  assign _T_443 = _T_245 ? 2'h0 : _T_442; // @[Lookup.scala 11:37:Sodor3Stage.fir@778.4]
  assign _T_444 = _T_241 ? 2'h2 : _T_443; // @[Lookup.scala 11:37:Sodor3Stage.fir@779.4]
  assign _T_445 = _T_237 ? 2'h2 : _T_444; // @[Lookup.scala 11:37:Sodor3Stage.fir@780.4]
  assign _T_446 = _T_233 ? 2'h0 : _T_445; // @[Lookup.scala 11:37:Sodor3Stage.fir@781.4]
  assign _T_447 = _T_229 ? 2'h0 : _T_446; // @[Lookup.scala 11:37:Sodor3Stage.fir@782.4]
  assign _T_448 = _T_225 ? 2'h0 : _T_447; // @[Lookup.scala 11:37:Sodor3Stage.fir@783.4]
  assign _T_449 = _T_221 ? 2'h0 : _T_448; // @[Lookup.scala 11:37:Sodor3Stage.fir@784.4]
  assign _T_450 = _T_217 ? 2'h0 : _T_449; // @[Lookup.scala 11:37:Sodor3Stage.fir@785.4]
  assign _T_451 = _T_213 ? 2'h0 : _T_450; // @[Lookup.scala 11:37:Sodor3Stage.fir@786.4]
  assign _T_452 = _T_209 ? 2'h0 : _T_451; // @[Lookup.scala 11:37:Sodor3Stage.fir@787.4]
  assign _T_453 = _T_205 ? 2'h0 : _T_452; // @[Lookup.scala 11:37:Sodor3Stage.fir@788.4]
  assign _T_454 = _T_201 ? 2'h0 : _T_453; // @[Lookup.scala 11:37:Sodor3Stage.fir@789.4]
  assign _T_455 = _T_197 ? 2'h0 : _T_454; // @[Lookup.scala 11:37:Sodor3Stage.fir@790.4]
  assign _T_456 = _T_193 ? 2'h0 : _T_455; // @[Lookup.scala 11:37:Sodor3Stage.fir@791.4]
  assign _T_457 = _T_189 ? 2'h0 : _T_456; // @[Lookup.scala 11:37:Sodor3Stage.fir@792.4]
  assign _T_458 = _T_185 ? 2'h0 : _T_457; // @[Lookup.scala 11:37:Sodor3Stage.fir@793.4]
  assign _T_459 = _T_181 ? 2'h0 : _T_458; // @[Lookup.scala 11:37:Sodor3Stage.fir@794.4]
  assign _T_460 = _T_177 ? 2'h0 : _T_459; // @[Lookup.scala 11:37:Sodor3Stage.fir@795.4]
  assign _T_461 = _T_173 ? 2'h0 : _T_460; // @[Lookup.scala 11:37:Sodor3Stage.fir@796.4]
  assign _T_462 = _T_169 ? 2'h0 : _T_461; // @[Lookup.scala 11:37:Sodor3Stage.fir@797.4]
  assign _T_463 = _T_165 ? 2'h0 : _T_462; // @[Lookup.scala 11:37:Sodor3Stage.fir@798.4]
  assign _T_464 = _T_161 ? 2'h0 : _T_463; // @[Lookup.scala 11:37:Sodor3Stage.fir@799.4]
  assign _T_465 = _T_157 ? 2'h0 : _T_464; // @[Lookup.scala 11:37:Sodor3Stage.fir@800.4]
  assign _T_466 = _T_153 ? 2'h0 : _T_465; // @[Lookup.scala 11:37:Sodor3Stage.fir@801.4]
  assign _T_467 = _T_149 ? 2'h0 : _T_466; // @[Lookup.scala 11:37:Sodor3Stage.fir@802.4]
  assign _T_468 = _T_145 ? 2'h0 : _T_467; // @[Lookup.scala 11:37:Sodor3Stage.fir@803.4]
  assign _T_469 = _T_141 ? 2'h0 : _T_468; // @[Lookup.scala 11:37:Sodor3Stage.fir@804.4]
  assign _T_470 = _T_137 ? 2'h0 : _T_469; // @[Lookup.scala 11:37:Sodor3Stage.fir@805.4]
  assign _T_471 = _T_133 ? 2'h0 : _T_470; // @[Lookup.scala 11:37:Sodor3Stage.fir@806.4]
  assign _T_472 = _T_129 ? 2'h0 : _T_471; // @[Lookup.scala 11:37:Sodor3Stage.fir@807.4]
  assign _T_473 = _T_125 ? 2'h1 : _T_472; // @[Lookup.scala 11:37:Sodor3Stage.fir@808.4]
  assign _T_474 = _T_121 ? 2'h1 : _T_473; // @[Lookup.scala 11:37:Sodor3Stage.fir@809.4]
  assign _T_475 = _T_117 ? 2'h0 : _T_474; // @[Lookup.scala 11:37:Sodor3Stage.fir@810.4]
  assign _T_476 = _T_113 ? 2'h0 : _T_475; // @[Lookup.scala 11:37:Sodor3Stage.fir@811.4]
  assign _T_477 = _T_109 ? 2'h0 : _T_476; // @[Lookup.scala 11:37:Sodor3Stage.fir@812.4]
  assign _T_478 = _T_105 ? 2'h0 : _T_477; // @[Lookup.scala 11:37:Sodor3Stage.fir@813.4]
  assign _T_479 = _T_101 ? 2'h0 : _T_478; // @[Lookup.scala 11:37:Sodor3Stage.fir@814.4]
  assign _T_480 = _T_97 ? 2'h0 : _T_479; // @[Lookup.scala 11:37:Sodor3Stage.fir@815.4]
  assign _T_481 = _T_93 ? 2'h0 : _T_480; // @[Lookup.scala 11:37:Sodor3Stage.fir@816.4]
  assign _T_501 = _T_209 ? 2'h1 : 2'h0; // @[Lookup.scala 11:37:Sodor3Stage.fir@837.4]
  assign _T_502 = _T_205 ? 2'h0 : _T_501; // @[Lookup.scala 11:37:Sodor3Stage.fir@838.4]
  assign _T_503 = _T_201 ? 2'h0 : _T_502; // @[Lookup.scala 11:37:Sodor3Stage.fir@839.4]
  assign _T_504 = _T_197 ? 2'h0 : _T_503; // @[Lookup.scala 11:37:Sodor3Stage.fir@840.4]
  assign _T_505 = _T_193 ? 2'h0 : _T_504; // @[Lookup.scala 11:37:Sodor3Stage.fir@841.4]
  assign _T_506 = _T_189 ? 2'h0 : _T_505; // @[Lookup.scala 11:37:Sodor3Stage.fir@842.4]
  assign _T_507 = _T_185 ? 2'h0 : _T_506; // @[Lookup.scala 11:37:Sodor3Stage.fir@843.4]
  assign _T_508 = _T_181 ? 2'h0 : _T_507; // @[Lookup.scala 11:37:Sodor3Stage.fir@844.4]
  assign _T_509 = _T_177 ? 2'h0 : _T_508; // @[Lookup.scala 11:37:Sodor3Stage.fir@845.4]
  assign _T_510 = _T_173 ? 2'h0 : _T_509; // @[Lookup.scala 11:37:Sodor3Stage.fir@846.4]
  assign _T_511 = _T_169 ? 2'h0 : _T_510; // @[Lookup.scala 11:37:Sodor3Stage.fir@847.4]
  assign _T_512 = _T_165 ? 2'h0 : _T_511; // @[Lookup.scala 11:37:Sodor3Stage.fir@848.4]
  assign _T_513 = _T_161 ? 2'h1 : _T_512; // @[Lookup.scala 11:37:Sodor3Stage.fir@849.4]
  assign _T_514 = _T_157 ? 2'h1 : _T_513; // @[Lookup.scala 11:37:Sodor3Stage.fir@850.4]
  assign _T_515 = _T_153 ? 2'h1 : _T_514; // @[Lookup.scala 11:37:Sodor3Stage.fir@851.4]
  assign _T_516 = _T_149 ? 2'h1 : _T_515; // @[Lookup.scala 11:37:Sodor3Stage.fir@852.4]
  assign _T_517 = _T_145 ? 2'h1 : _T_516; // @[Lookup.scala 11:37:Sodor3Stage.fir@853.4]
  assign _T_518 = _T_141 ? 2'h1 : _T_517; // @[Lookup.scala 11:37:Sodor3Stage.fir@854.4]
  assign _T_519 = _T_137 ? 2'h1 : _T_518; // @[Lookup.scala 11:37:Sodor3Stage.fir@855.4]
  assign _T_520 = _T_133 ? 2'h1 : _T_519; // @[Lookup.scala 11:37:Sodor3Stage.fir@856.4]
  assign _T_521 = _T_129 ? 2'h1 : _T_520; // @[Lookup.scala 11:37:Sodor3Stage.fir@857.4]
  assign _T_522 = _T_125 ? 2'h0 : _T_521; // @[Lookup.scala 11:37:Sodor3Stage.fir@858.4]
  assign _T_523 = _T_121 ? 2'h3 : _T_522; // @[Lookup.scala 11:37:Sodor3Stage.fir@859.4]
  assign _T_524 = _T_117 ? 2'h2 : _T_523; // @[Lookup.scala 11:37:Sodor3Stage.fir@860.4]
  assign _T_525 = _T_113 ? 2'h2 : _T_524; // @[Lookup.scala 11:37:Sodor3Stage.fir@861.4]
  assign _T_526 = _T_109 ? 2'h2 : _T_525; // @[Lookup.scala 11:37:Sodor3Stage.fir@862.4]
  assign _T_527 = _T_105 ? 2'h1 : _T_526; // @[Lookup.scala 11:37:Sodor3Stage.fir@863.4]
  assign _T_528 = _T_101 ? 2'h1 : _T_527; // @[Lookup.scala 11:37:Sodor3Stage.fir@864.4]
  assign _T_529 = _T_97 ? 2'h1 : _T_528; // @[Lookup.scala 11:37:Sodor3Stage.fir@865.4]
  assign _T_530 = _T_93 ? 2'h1 : _T_529; // @[Lookup.scala 11:37:Sodor3Stage.fir@866.4]
  assign _T_538 = _T_257 ? 4'h8 : 4'h0; // @[Lookup.scala 11:37:Sodor3Stage.fir@875.4]
  assign _T_539 = _T_253 ? 4'h8 : _T_538; // @[Lookup.scala 11:37:Sodor3Stage.fir@876.4]
  assign _T_540 = _T_249 ? 4'h8 : _T_539; // @[Lookup.scala 11:37:Sodor3Stage.fir@877.4]
  assign _T_541 = _T_245 ? 4'h8 : _T_540; // @[Lookup.scala 11:37:Sodor3Stage.fir@878.4]
  assign _T_542 = _T_241 ? 4'h8 : _T_541; // @[Lookup.scala 11:37:Sodor3Stage.fir@879.4]
  assign _T_543 = _T_237 ? 4'h8 : _T_542; // @[Lookup.scala 11:37:Sodor3Stage.fir@880.4]
  assign _T_544 = _T_233 ? 4'h0 : _T_543; // @[Lookup.scala 11:37:Sodor3Stage.fir@881.4]
  assign _T_545 = _T_229 ? 4'h0 : _T_544; // @[Lookup.scala 11:37:Sodor3Stage.fir@882.4]
  assign _T_546 = _T_225 ? 4'h0 : _T_545; // @[Lookup.scala 11:37:Sodor3Stage.fir@883.4]
  assign _T_547 = _T_221 ? 4'h0 : _T_546; // @[Lookup.scala 11:37:Sodor3Stage.fir@884.4]
  assign _T_548 = _T_217 ? 4'h0 : _T_547; // @[Lookup.scala 11:37:Sodor3Stage.fir@885.4]
  assign _T_549 = _T_213 ? 4'h0 : _T_548; // @[Lookup.scala 11:37:Sodor3Stage.fir@886.4]
  assign _T_550 = _T_209 ? 4'h0 : _T_549; // @[Lookup.scala 11:37:Sodor3Stage.fir@887.4]
  assign _T_551 = _T_205 ? 4'h0 : _T_550; // @[Lookup.scala 11:37:Sodor3Stage.fir@888.4]
  assign _T_552 = _T_201 ? 4'h5 : _T_551; // @[Lookup.scala 11:37:Sodor3Stage.fir@889.4]
  assign _T_553 = _T_197 ? 4'hb : _T_552; // @[Lookup.scala 11:37:Sodor3Stage.fir@890.4]
  assign _T_554 = _T_193 ? 4'h4 : _T_553; // @[Lookup.scala 11:37:Sodor3Stage.fir@891.4]
  assign _T_555 = _T_189 ? 4'h6 : _T_554; // @[Lookup.scala 11:37:Sodor3Stage.fir@892.4]
  assign _T_556 = _T_185 ? 4'h7 : _T_555; // @[Lookup.scala 11:37:Sodor3Stage.fir@893.4]
  assign _T_557 = _T_181 ? 4'he : _T_556; // @[Lookup.scala 11:37:Sodor3Stage.fir@894.4]
  assign _T_558 = _T_177 ? 4'hc : _T_557; // @[Lookup.scala 11:37:Sodor3Stage.fir@895.4]
  assign _T_559 = _T_173 ? 4'ha : _T_558; // @[Lookup.scala 11:37:Sodor3Stage.fir@896.4]
  assign _T_560 = _T_169 ? 4'h0 : _T_559; // @[Lookup.scala 11:37:Sodor3Stage.fir@897.4]
  assign _T_561 = _T_165 ? 4'h1 : _T_560; // @[Lookup.scala 11:37:Sodor3Stage.fir@898.4]
  assign _T_562 = _T_161 ? 4'h5 : _T_561; // @[Lookup.scala 11:37:Sodor3Stage.fir@899.4]
  assign _T_563 = _T_157 ? 4'hb : _T_562; // @[Lookup.scala 11:37:Sodor3Stage.fir@900.4]
  assign _T_564 = _T_153 ? 4'h1 : _T_563; // @[Lookup.scala 11:37:Sodor3Stage.fir@901.4]
  assign _T_565 = _T_149 ? 4'he : _T_564; // @[Lookup.scala 11:37:Sodor3Stage.fir@902.4]
  assign _T_566 = _T_145 ? 4'hc : _T_565; // @[Lookup.scala 11:37:Sodor3Stage.fir@903.4]
  assign _T_567 = _T_141 ? 4'h4 : _T_566; // @[Lookup.scala 11:37:Sodor3Stage.fir@904.4]
  assign _T_568 = _T_137 ? 4'h6 : _T_567; // @[Lookup.scala 11:37:Sodor3Stage.fir@905.4]
  assign _T_569 = _T_133 ? 4'h7 : _T_568; // @[Lookup.scala 11:37:Sodor3Stage.fir@906.4]
  assign _T_570 = _T_129 ? 4'h0 : _T_569; // @[Lookup.scala 11:37:Sodor3Stage.fir@907.4]
  assign _T_571 = _T_125 ? 4'h8 : _T_570; // @[Lookup.scala 11:37:Sodor3Stage.fir@908.4]
  assign _T_572 = _T_121 ? 4'h0 : _T_571; // @[Lookup.scala 11:37:Sodor3Stage.fir@909.4]
  assign _T_573 = _T_117 ? 4'h0 : _T_572; // @[Lookup.scala 11:37:Sodor3Stage.fir@910.4]
  assign _T_574 = _T_113 ? 4'h0 : _T_573; // @[Lookup.scala 11:37:Sodor3Stage.fir@911.4]
  assign _T_575 = _T_109 ? 4'h0 : _T_574; // @[Lookup.scala 11:37:Sodor3Stage.fir@912.4]
  assign _T_576 = _T_105 ? 4'h0 : _T_575; // @[Lookup.scala 11:37:Sodor3Stage.fir@913.4]
  assign _T_577 = _T_101 ? 4'h0 : _T_576; // @[Lookup.scala 11:37:Sodor3Stage.fir@914.4]
  assign _T_578 = _T_97 ? 4'h0 : _T_577; // @[Lookup.scala 11:37:Sodor3Stage.fir@915.4]
  assign _T_579 = _T_93 ? 4'h0 : _T_578; // @[Lookup.scala 11:37:Sodor3Stage.fir@916.4]
  assign _T_587 = _T_257 ? 2'h3 : 2'h0; // @[Lookup.scala 11:37:Sodor3Stage.fir@925.4]
  assign _T_588 = _T_253 ? 2'h3 : _T_587; // @[Lookup.scala 11:37:Sodor3Stage.fir@926.4]
  assign _T_589 = _T_249 ? 2'h3 : _T_588; // @[Lookup.scala 11:37:Sodor3Stage.fir@927.4]
  assign _T_590 = _T_245 ? 2'h3 : _T_589; // @[Lookup.scala 11:37:Sodor3Stage.fir@928.4]
  assign _T_591 = _T_241 ? 2'h3 : _T_590; // @[Lookup.scala 11:37:Sodor3Stage.fir@929.4]
  assign _T_592 = _T_237 ? 2'h3 : _T_591; // @[Lookup.scala 11:37:Sodor3Stage.fir@930.4]
  assign _T_593 = _T_233 ? 2'h0 : _T_592; // @[Lookup.scala 11:37:Sodor3Stage.fir@931.4]
  assign _T_594 = _T_229 ? 2'h0 : _T_593; // @[Lookup.scala 11:37:Sodor3Stage.fir@932.4]
  assign _T_595 = _T_225 ? 2'h0 : _T_594; // @[Lookup.scala 11:37:Sodor3Stage.fir@933.4]
  assign _T_596 = _T_221 ? 2'h0 : _T_595; // @[Lookup.scala 11:37:Sodor3Stage.fir@934.4]
  assign _T_597 = _T_217 ? 2'h0 : _T_596; // @[Lookup.scala 11:37:Sodor3Stage.fir@935.4]
  assign _T_598 = _T_213 ? 2'h0 : _T_597; // @[Lookup.scala 11:37:Sodor3Stage.fir@936.4]
  assign _T_599 = _T_209 ? 2'h2 : _T_598; // @[Lookup.scala 11:37:Sodor3Stage.fir@937.4]
  assign _T_600 = _T_205 ? 2'h2 : _T_599; // @[Lookup.scala 11:37:Sodor3Stage.fir@938.4]
  assign _T_601 = _T_201 ? 2'h0 : _T_600; // @[Lookup.scala 11:37:Sodor3Stage.fir@939.4]
  assign _T_602 = _T_197 ? 2'h0 : _T_601; // @[Lookup.scala 11:37:Sodor3Stage.fir@940.4]
  assign _T_603 = _T_193 ? 2'h0 : _T_602; // @[Lookup.scala 11:37:Sodor3Stage.fir@941.4]
  assign _T_604 = _T_189 ? 2'h0 : _T_603; // @[Lookup.scala 11:37:Sodor3Stage.fir@942.4]
  assign _T_605 = _T_185 ? 2'h0 : _T_604; // @[Lookup.scala 11:37:Sodor3Stage.fir@943.4]
  assign _T_606 = _T_181 ? 2'h0 : _T_605; // @[Lookup.scala 11:37:Sodor3Stage.fir@944.4]
  assign _T_607 = _T_177 ? 2'h0 : _T_606; // @[Lookup.scala 11:37:Sodor3Stage.fir@945.4]
  assign _T_608 = _T_173 ? 2'h0 : _T_607; // @[Lookup.scala 11:37:Sodor3Stage.fir@946.4]
  assign _T_609 = _T_169 ? 2'h0 : _T_608; // @[Lookup.scala 11:37:Sodor3Stage.fir@947.4]
  assign _T_610 = _T_165 ? 2'h0 : _T_609; // @[Lookup.scala 11:37:Sodor3Stage.fir@948.4]
  assign _T_611 = _T_161 ? 2'h0 : _T_610; // @[Lookup.scala 11:37:Sodor3Stage.fir@949.4]
  assign _T_612 = _T_157 ? 2'h0 : _T_611; // @[Lookup.scala 11:37:Sodor3Stage.fir@950.4]
  assign _T_613 = _T_153 ? 2'h0 : _T_612; // @[Lookup.scala 11:37:Sodor3Stage.fir@951.4]
  assign _T_614 = _T_149 ? 2'h0 : _T_613; // @[Lookup.scala 11:37:Sodor3Stage.fir@952.4]
  assign _T_615 = _T_145 ? 2'h0 : _T_614; // @[Lookup.scala 11:37:Sodor3Stage.fir@953.4]
  assign _T_616 = _T_141 ? 2'h0 : _T_615; // @[Lookup.scala 11:37:Sodor3Stage.fir@954.4]
  assign _T_617 = _T_137 ? 2'h0 : _T_616; // @[Lookup.scala 11:37:Sodor3Stage.fir@955.4]
  assign _T_618 = _T_133 ? 2'h0 : _T_617; // @[Lookup.scala 11:37:Sodor3Stage.fir@956.4]
  assign _T_619 = _T_129 ? 2'h0 : _T_618; // @[Lookup.scala 11:37:Sodor3Stage.fir@957.4]
  assign _T_620 = _T_125 ? 2'h0 : _T_619; // @[Lookup.scala 11:37:Sodor3Stage.fir@958.4]
  assign _T_621 = _T_121 ? 2'h0 : _T_620; // @[Lookup.scala 11:37:Sodor3Stage.fir@959.4]
  assign _T_622 = _T_117 ? 2'h0 : _T_621; // @[Lookup.scala 11:37:Sodor3Stage.fir@960.4]
  assign _T_623 = _T_113 ? 2'h0 : _T_622; // @[Lookup.scala 11:37:Sodor3Stage.fir@961.4]
  assign _T_624 = _T_109 ? 2'h0 : _T_623; // @[Lookup.scala 11:37:Sodor3Stage.fir@962.4]
  assign _T_625 = _T_105 ? 2'h1 : _T_624; // @[Lookup.scala 11:37:Sodor3Stage.fir@963.4]
  assign _T_626 = _T_101 ? 2'h1 : _T_625; // @[Lookup.scala 11:37:Sodor3Stage.fir@964.4]
  assign _T_627 = _T_97 ? 2'h1 : _T_626; // @[Lookup.scala 11:37:Sodor3Stage.fir@965.4]
  assign _T_628 = _T_93 ? 2'h1 : _T_627; // @[Lookup.scala 11:37:Sodor3Stage.fir@966.4]
  assign _T_637 = _T_253 ? 1'h1 : _T_257; // @[Lookup.scala 11:37:Sodor3Stage.fir@976.4]
  assign _T_638 = _T_249 ? 1'h1 : _T_637; // @[Lookup.scala 11:37:Sodor3Stage.fir@977.4]
  assign _T_639 = _T_245 ? 1'h1 : _T_638; // @[Lookup.scala 11:37:Sodor3Stage.fir@978.4]
  assign _T_640 = _T_241 ? 1'h1 : _T_639; // @[Lookup.scala 11:37:Sodor3Stage.fir@979.4]
  assign _T_641 = _T_237 ? 1'h1 : _T_640; // @[Lookup.scala 11:37:Sodor3Stage.fir@980.4]
  assign _T_642 = _T_233 ? 1'h0 : _T_641; // @[Lookup.scala 11:37:Sodor3Stage.fir@981.4]
  assign _T_643 = _T_229 ? 1'h0 : _T_642; // @[Lookup.scala 11:37:Sodor3Stage.fir@982.4]
  assign _T_644 = _T_225 ? 1'h0 : _T_643; // @[Lookup.scala 11:37:Sodor3Stage.fir@983.4]
  assign _T_645 = _T_221 ? 1'h0 : _T_644; // @[Lookup.scala 11:37:Sodor3Stage.fir@984.4]
  assign _T_646 = _T_217 ? 1'h0 : _T_645; // @[Lookup.scala 11:37:Sodor3Stage.fir@985.4]
  assign _T_647 = _T_213 ? 1'h0 : _T_646; // @[Lookup.scala 11:37:Sodor3Stage.fir@986.4]
  assign _T_648 = _T_209 ? 1'h1 : _T_647; // @[Lookup.scala 11:37:Sodor3Stage.fir@987.4]
  assign _T_649 = _T_205 ? 1'h1 : _T_648; // @[Lookup.scala 11:37:Sodor3Stage.fir@988.4]
  assign _T_650 = _T_201 ? 1'h1 : _T_649; // @[Lookup.scala 11:37:Sodor3Stage.fir@989.4]
  assign _T_651 = _T_197 ? 1'h1 : _T_650; // @[Lookup.scala 11:37:Sodor3Stage.fir@990.4]
  assign _T_652 = _T_193 ? 1'h1 : _T_651; // @[Lookup.scala 11:37:Sodor3Stage.fir@991.4]
  assign _T_653 = _T_189 ? 1'h1 : _T_652; // @[Lookup.scala 11:37:Sodor3Stage.fir@992.4]
  assign _T_654 = _T_185 ? 1'h1 : _T_653; // @[Lookup.scala 11:37:Sodor3Stage.fir@993.4]
  assign _T_655 = _T_181 ? 1'h1 : _T_654; // @[Lookup.scala 11:37:Sodor3Stage.fir@994.4]
  assign _T_656 = _T_177 ? 1'h1 : _T_655; // @[Lookup.scala 11:37:Sodor3Stage.fir@995.4]
  assign _T_657 = _T_173 ? 1'h1 : _T_656; // @[Lookup.scala 11:37:Sodor3Stage.fir@996.4]
  assign _T_658 = _T_169 ? 1'h1 : _T_657; // @[Lookup.scala 11:37:Sodor3Stage.fir@997.4]
  assign _T_659 = _T_165 ? 1'h1 : _T_658; // @[Lookup.scala 11:37:Sodor3Stage.fir@998.4]
  assign _T_660 = _T_161 ? 1'h1 : _T_659; // @[Lookup.scala 11:37:Sodor3Stage.fir@999.4]
  assign _T_661 = _T_157 ? 1'h1 : _T_660; // @[Lookup.scala 11:37:Sodor3Stage.fir@1000.4]
  assign _T_662 = _T_153 ? 1'h1 : _T_661; // @[Lookup.scala 11:37:Sodor3Stage.fir@1001.4]
  assign _T_663 = _T_149 ? 1'h1 : _T_662; // @[Lookup.scala 11:37:Sodor3Stage.fir@1002.4]
  assign _T_664 = _T_145 ? 1'h1 : _T_663; // @[Lookup.scala 11:37:Sodor3Stage.fir@1003.4]
  assign _T_665 = _T_141 ? 1'h1 : _T_664; // @[Lookup.scala 11:37:Sodor3Stage.fir@1004.4]
  assign _T_666 = _T_137 ? 1'h1 : _T_665; // @[Lookup.scala 11:37:Sodor3Stage.fir@1005.4]
  assign _T_667 = _T_133 ? 1'h1 : _T_666; // @[Lookup.scala 11:37:Sodor3Stage.fir@1006.4]
  assign _T_668 = _T_129 ? 1'h1 : _T_667; // @[Lookup.scala 11:37:Sodor3Stage.fir@1007.4]
  assign _T_669 = _T_125 ? 1'h1 : _T_668; // @[Lookup.scala 11:37:Sodor3Stage.fir@1008.4]
  assign _T_670 = _T_121 ? 1'h1 : _T_669; // @[Lookup.scala 11:37:Sodor3Stage.fir@1009.4]
  assign _T_671 = _T_117 ? 1'h0 : _T_670; // @[Lookup.scala 11:37:Sodor3Stage.fir@1010.4]
  assign _T_672 = _T_113 ? 1'h0 : _T_671; // @[Lookup.scala 11:37:Sodor3Stage.fir@1011.4]
  assign _T_673 = _T_109 ? 1'h0 : _T_672; // @[Lookup.scala 11:37:Sodor3Stage.fir@1012.4]
  assign _T_674 = _T_105 ? 1'h1 : _T_673; // @[Lookup.scala 11:37:Sodor3Stage.fir@1013.4]
  assign _T_675 = _T_101 ? 1'h1 : _T_674; // @[Lookup.scala 11:37:Sodor3Stage.fir@1014.4]
  assign _T_676 = _T_97 ? 1'h1 : _T_675; // @[Lookup.scala 11:37:Sodor3Stage.fir@1015.4]
  assign _T_677 = _T_93 ? 1'h1 : _T_676; // @[Lookup.scala 11:37:Sodor3Stage.fir@1016.4]
  assign cs0_2 = _T_89 ? 1'h1 : _T_677; // @[Lookup.scala 11:37:Sodor3Stage.fir@1017.4]
  assign _T_699 = _T_201 ? 1'h1 : _T_205; // @[Lookup.scala 11:37:Sodor3Stage.fir@1039.4]
  assign _T_700 = _T_197 ? 1'h1 : _T_699; // @[Lookup.scala 11:37:Sodor3Stage.fir@1040.4]
  assign _T_701 = _T_193 ? 1'h1 : _T_700; // @[Lookup.scala 11:37:Sodor3Stage.fir@1041.4]
  assign _T_702 = _T_189 ? 1'h1 : _T_701; // @[Lookup.scala 11:37:Sodor3Stage.fir@1042.4]
  assign _T_703 = _T_185 ? 1'h1 : _T_702; // @[Lookup.scala 11:37:Sodor3Stage.fir@1043.4]
  assign _T_704 = _T_181 ? 1'h1 : _T_703; // @[Lookup.scala 11:37:Sodor3Stage.fir@1044.4]
  assign _T_705 = _T_177 ? 1'h1 : _T_704; // @[Lookup.scala 11:37:Sodor3Stage.fir@1045.4]
  assign _T_706 = _T_173 ? 1'h1 : _T_705; // @[Lookup.scala 11:37:Sodor3Stage.fir@1046.4]
  assign _T_707 = _T_169 ? 1'h1 : _T_706; // @[Lookup.scala 11:37:Sodor3Stage.fir@1047.4]
  assign _T_708 = _T_165 ? 1'h1 : _T_707; // @[Lookup.scala 11:37:Sodor3Stage.fir@1048.4]
  assign _T_709 = _T_161 ? 1'h1 : _T_708; // @[Lookup.scala 11:37:Sodor3Stage.fir@1049.4]
  assign _T_710 = _T_157 ? 1'h1 : _T_709; // @[Lookup.scala 11:37:Sodor3Stage.fir@1050.4]
  assign _T_711 = _T_153 ? 1'h1 : _T_710; // @[Lookup.scala 11:37:Sodor3Stage.fir@1051.4]
  assign _T_712 = _T_149 ? 1'h1 : _T_711; // @[Lookup.scala 11:37:Sodor3Stage.fir@1052.4]
  assign _T_713 = _T_145 ? 1'h1 : _T_712; // @[Lookup.scala 11:37:Sodor3Stage.fir@1053.4]
  assign _T_714 = _T_141 ? 1'h1 : _T_713; // @[Lookup.scala 11:37:Sodor3Stage.fir@1054.4]
  assign _T_715 = _T_137 ? 1'h1 : _T_714; // @[Lookup.scala 11:37:Sodor3Stage.fir@1055.4]
  assign _T_716 = _T_133 ? 1'h1 : _T_715; // @[Lookup.scala 11:37:Sodor3Stage.fir@1056.4]
  assign _T_717 = _T_129 ? 1'h1 : _T_716; // @[Lookup.scala 11:37:Sodor3Stage.fir@1057.4]
  assign _T_718 = _T_125 ? 1'h1 : _T_717; // @[Lookup.scala 11:37:Sodor3Stage.fir@1058.4]
  assign _T_719 = _T_121 ? 1'h1 : _T_718; // @[Lookup.scala 11:37:Sodor3Stage.fir@1059.4]
  assign _T_720 = _T_117 ? 1'h0 : _T_719; // @[Lookup.scala 11:37:Sodor3Stage.fir@1060.4]
  assign _T_721 = _T_113 ? 1'h0 : _T_720; // @[Lookup.scala 11:37:Sodor3Stage.fir@1061.4]
  assign _T_722 = _T_109 ? 1'h0 : _T_721; // @[Lookup.scala 11:37:Sodor3Stage.fir@1062.4]
  assign _T_723 = _T_105 ? 1'h0 : _T_722; // @[Lookup.scala 11:37:Sodor3Stage.fir@1063.4]
  assign _T_724 = _T_101 ? 1'h0 : _T_723; // @[Lookup.scala 11:37:Sodor3Stage.fir@1064.4]
  assign _T_725 = _T_97 ? 1'h0 : _T_724; // @[Lookup.scala 11:37:Sodor3Stage.fir@1065.4]
  assign _T_726 = _T_93 ? 1'h0 : _T_725; // @[Lookup.scala 11:37:Sodor3Stage.fir@1066.4]
  assign _T_819 = _T_113 ? 1'h1 : _T_117; // @[Lookup.scala 11:37:Sodor3Stage.fir@1161.4]
  assign _T_820 = _T_109 ? 1'h1 : _T_819; // @[Lookup.scala 11:37:Sodor3Stage.fir@1162.4]
  assign _T_821 = _T_105 ? 1'h0 : _T_820; // @[Lookup.scala 11:37:Sodor3Stage.fir@1163.4]
  assign _T_822 = _T_101 ? 1'h0 : _T_821; // @[Lookup.scala 11:37:Sodor3Stage.fir@1164.4]
  assign _T_823 = _T_97 ? 1'h0 : _T_822; // @[Lookup.scala 11:37:Sodor3Stage.fir@1165.4]
  assign _T_824 = _T_93 ? 1'h0 : _T_823; // @[Lookup.scala 11:37:Sodor3Stage.fir@1166.4]
  assign _T_867 = _T_117 ? 3'h2 : 3'h0; // @[Lookup.scala 11:37:Sodor3Stage.fir@1210.4]
  assign _T_868 = _T_113 ? 3'h1 : _T_867; // @[Lookup.scala 11:37:Sodor3Stage.fir@1211.4]
  assign _T_869 = _T_109 ? 3'h3 : _T_868; // @[Lookup.scala 11:37:Sodor3Stage.fir@1212.4]
  assign _T_870 = _T_105 ? 3'h6 : _T_869; // @[Lookup.scala 11:37:Sodor3Stage.fir@1213.4]
  assign _T_871 = _T_101 ? 3'h2 : _T_870; // @[Lookup.scala 11:37:Sodor3Stage.fir@1214.4]
  assign _T_872 = _T_97 ? 3'h5 : _T_871; // @[Lookup.scala 11:37:Sodor3Stage.fir@1215.4]
  assign _T_873 = _T_93 ? 3'h1 : _T_872; // @[Lookup.scala 11:37:Sodor3Stage.fir@1216.4]
  assign _T_876 = _T_277 ? 3'h4 : 3'h0; // @[Lookup.scala 11:37:Sodor3Stage.fir@1220.4]
  assign _T_877 = _T_273 ? 3'h4 : _T_876; // @[Lookup.scala 11:37:Sodor3Stage.fir@1221.4]
  assign _T_878 = _T_269 ? 3'h4 : _T_877; // @[Lookup.scala 11:37:Sodor3Stage.fir@1222.4]
  assign _T_879 = _T_265 ? 3'h4 : _T_878; // @[Lookup.scala 11:37:Sodor3Stage.fir@1223.4]
  assign _T_880 = _T_261 ? 3'h4 : _T_879; // @[Lookup.scala 11:37:Sodor3Stage.fir@1224.4]
  assign _T_881 = _T_257 ? 3'h3 : _T_880; // @[Lookup.scala 11:37:Sodor3Stage.fir@1225.4]
  assign _T_882 = _T_253 ? 3'h3 : _T_881; // @[Lookup.scala 11:37:Sodor3Stage.fir@1226.4]
  assign _T_883 = _T_249 ? 3'h2 : _T_882; // @[Lookup.scala 11:37:Sodor3Stage.fir@1227.4]
  assign _T_884 = _T_245 ? 3'h1 : _T_883; // @[Lookup.scala 11:37:Sodor3Stage.fir@1228.4]
  assign _T_885 = _T_241 ? 3'h2 : _T_884; // @[Lookup.scala 11:37:Sodor3Stage.fir@1229.4]
  assign _T_886 = _T_237 ? 3'h1 : _T_885; // @[Lookup.scala 11:37:Sodor3Stage.fir@1230.4]
  assign _T_887 = _T_233 ? 3'h0 : _T_886; // @[Lookup.scala 11:37:Sodor3Stage.fir@1231.4]
  assign _T_888 = _T_229 ? 3'h0 : _T_887; // @[Lookup.scala 11:37:Sodor3Stage.fir@1232.4]
  assign _T_889 = _T_225 ? 3'h0 : _T_888; // @[Lookup.scala 11:37:Sodor3Stage.fir@1233.4]
  assign _T_890 = _T_221 ? 3'h0 : _T_889; // @[Lookup.scala 11:37:Sodor3Stage.fir@1234.4]
  assign _T_891 = _T_217 ? 3'h0 : _T_890; // @[Lookup.scala 11:37:Sodor3Stage.fir@1235.4]
  assign _T_892 = _T_213 ? 3'h0 : _T_891; // @[Lookup.scala 11:37:Sodor3Stage.fir@1236.4]
  assign _T_893 = _T_209 ? 3'h0 : _T_892; // @[Lookup.scala 11:37:Sodor3Stage.fir@1237.4]
  assign _T_894 = _T_205 ? 3'h0 : _T_893; // @[Lookup.scala 11:37:Sodor3Stage.fir@1238.4]
  assign _T_895 = _T_201 ? 3'h0 : _T_894; // @[Lookup.scala 11:37:Sodor3Stage.fir@1239.4]
  assign _T_896 = _T_197 ? 3'h0 : _T_895; // @[Lookup.scala 11:37:Sodor3Stage.fir@1240.4]
  assign _T_897 = _T_193 ? 3'h0 : _T_896; // @[Lookup.scala 11:37:Sodor3Stage.fir@1241.4]
  assign _T_898 = _T_189 ? 3'h0 : _T_897; // @[Lookup.scala 11:37:Sodor3Stage.fir@1242.4]
  assign _T_899 = _T_185 ? 3'h0 : _T_898; // @[Lookup.scala 11:37:Sodor3Stage.fir@1243.4]
  assign _T_900 = _T_181 ? 3'h0 : _T_899; // @[Lookup.scala 11:37:Sodor3Stage.fir@1244.4]
  assign _T_901 = _T_177 ? 3'h0 : _T_900; // @[Lookup.scala 11:37:Sodor3Stage.fir@1245.4]
  assign _T_902 = _T_173 ? 3'h0 : _T_901; // @[Lookup.scala 11:37:Sodor3Stage.fir@1246.4]
  assign _T_903 = _T_169 ? 3'h0 : _T_902; // @[Lookup.scala 11:37:Sodor3Stage.fir@1247.4]
  assign _T_904 = _T_165 ? 3'h0 : _T_903; // @[Lookup.scala 11:37:Sodor3Stage.fir@1248.4]
  assign _T_905 = _T_161 ? 3'h0 : _T_904; // @[Lookup.scala 11:37:Sodor3Stage.fir@1249.4]
  assign _T_906 = _T_157 ? 3'h0 : _T_905; // @[Lookup.scala 11:37:Sodor3Stage.fir@1250.4]
  assign _T_907 = _T_153 ? 3'h0 : _T_906; // @[Lookup.scala 11:37:Sodor3Stage.fir@1251.4]
  assign _T_908 = _T_149 ? 3'h0 : _T_907; // @[Lookup.scala 11:37:Sodor3Stage.fir@1252.4]
  assign _T_909 = _T_145 ? 3'h0 : _T_908; // @[Lookup.scala 11:37:Sodor3Stage.fir@1253.4]
  assign _T_910 = _T_141 ? 3'h0 : _T_909; // @[Lookup.scala 11:37:Sodor3Stage.fir@1254.4]
  assign _T_911 = _T_137 ? 3'h0 : _T_910; // @[Lookup.scala 11:37:Sodor3Stage.fir@1255.4]
  assign _T_912 = _T_133 ? 3'h0 : _T_911; // @[Lookup.scala 11:37:Sodor3Stage.fir@1256.4]
  assign _T_913 = _T_129 ? 3'h0 : _T_912; // @[Lookup.scala 11:37:Sodor3Stage.fir@1257.4]
  assign _T_914 = _T_125 ? 3'h0 : _T_913; // @[Lookup.scala 11:37:Sodor3Stage.fir@1258.4]
  assign _T_915 = _T_121 ? 3'h0 : _T_914; // @[Lookup.scala 11:37:Sodor3Stage.fir@1259.4]
  assign _T_916 = _T_117 ? 3'h0 : _T_915; // @[Lookup.scala 11:37:Sodor3Stage.fir@1260.4]
  assign _T_917 = _T_113 ? 3'h0 : _T_916; // @[Lookup.scala 11:37:Sodor3Stage.fir@1261.4]
  assign _T_918 = _T_109 ? 3'h0 : _T_917; // @[Lookup.scala 11:37:Sodor3Stage.fir@1262.4]
  assign _T_919 = _T_105 ? 3'h0 : _T_918; // @[Lookup.scala 11:37:Sodor3Stage.fir@1263.4]
  assign _T_920 = _T_101 ? 3'h0 : _T_919; // @[Lookup.scala 11:37:Sodor3Stage.fir@1264.4]
  assign _T_921 = _T_97 ? 3'h0 : _T_920; // @[Lookup.scala 11:37:Sodor3Stage.fir@1265.4]
  assign _T_922 = _T_93 ? 3'h0 : _T_921; // @[Lookup.scala 11:37:Sodor3Stage.fir@1266.4]
  assign cs0_7 = _T_89 ? 3'h0 : _T_922; // @[Lookup.scala 11:37:Sodor3Stage.fir@1267.4]
  assign _T_973 = cs_br_type == 4'h0; // @[cpath.scala 138:37:Sodor3Stage.fir@1319.4]
  assign _T_974 = cs_br_type == 4'h1; // @[cpath.scala 139:37:Sodor3Stage.fir@1320.4]
  assign _T_976 = io_dat_br_eq == 1'h0; // @[cpath.scala 139:54:Sodor3Stage.fir@1321.4]
  assign _T_977 = _T_976 ? 3'h1 : 3'h0; // @[cpath.scala 139:53:Sodor3Stage.fir@1322.4]
  assign _T_978 = cs_br_type == 4'h2; // @[cpath.scala 140:37:Sodor3Stage.fir@1323.4]
  assign _T_979 = io_dat_br_eq ? 3'h1 : 3'h0; // @[cpath.scala 140:53:Sodor3Stage.fir@1324.4]
  assign _T_980 = cs_br_type == 4'h3; // @[cpath.scala 141:37:Sodor3Stage.fir@1325.4]
  assign _T_982 = io_dat_br_lt == 1'h0; // @[cpath.scala 141:54:Sodor3Stage.fir@1326.4]
  assign _T_983 = _T_982 ? 3'h1 : 3'h0; // @[cpath.scala 141:53:Sodor3Stage.fir@1327.4]
  assign _T_984 = cs_br_type == 4'h4; // @[cpath.scala 142:37:Sodor3Stage.fir@1328.4]
  assign _T_986 = io_dat_br_ltu == 1'h0; // @[cpath.scala 142:54:Sodor3Stage.fir@1329.4]
  assign _T_987 = _T_986 ? 3'h1 : 3'h0; // @[cpath.scala 142:53:Sodor3Stage.fir@1330.4]
  assign _T_988 = cs_br_type == 4'h5; // @[cpath.scala 143:37:Sodor3Stage.fir@1331.4]
  assign _T_989 = io_dat_br_lt ? 3'h1 : 3'h0; // @[cpath.scala 143:53:Sodor3Stage.fir@1332.4]
  assign _T_990 = cs_br_type == 4'h6; // @[cpath.scala 144:37:Sodor3Stage.fir@1333.4]
  assign _T_991 = io_dat_br_ltu ? 3'h1 : 3'h0; // @[cpath.scala 144:53:Sodor3Stage.fir@1334.4]
  assign _T_992 = cs_br_type == 4'h7; // @[cpath.scala 145:37:Sodor3Stage.fir@1335.4]
  assign _T_993 = cs_br_type == 4'h8; // @[cpath.scala 146:37:Sodor3Stage.fir@1336.4]
  assign _T_994 = _T_993 ? 3'h3 : 3'h0; // @[cpath.scala 146:25:Sodor3Stage.fir@1337.4]
  assign _T_995 = _T_992 ? 3'h2 : _T_994; // @[cpath.scala 145:25:Sodor3Stage.fir@1338.4]
  assign _T_996 = _T_990 ? _T_991 : _T_995; // @[cpath.scala 144:25:Sodor3Stage.fir@1339.4]
  assign _T_997 = _T_988 ? _T_989 : _T_996; // @[cpath.scala 143:25:Sodor3Stage.fir@1340.4]
  assign _T_998 = _T_984 ? _T_987 : _T_997; // @[cpath.scala 142:25:Sodor3Stage.fir@1341.4]
  assign _T_999 = _T_980 ? _T_983 : _T_998; // @[cpath.scala 141:25:Sodor3Stage.fir@1342.4]
  assign _T_1000 = _T_978 ? _T_979 : _T_999; // @[cpath.scala 140:25:Sodor3Stage.fir@1343.4]
  assign _T_1001 = _T_974 ? _T_977 : _T_1000; // @[cpath.scala 139:25:Sodor3Stage.fir@1344.4]
  assign _T_1002 = _T_973 ? 3'h0 : _T_1001; // @[cpath.scala 138:25:Sodor3Stage.fir@1345.4]
  assign take_evec = _T_1028 | io_dat_csr_eret; // @[cpath.scala 179:51:Sodor3Stage.fir@1385.4]
  assign ctrl_pc_sel = take_evec ? 3'h4 : _T_1002; // @[cpath.scala 137:25:Sodor3Stage.fir@1346.4]
  assign _T_1003 = ctrl_pc_sel == 3'h0; // @[cpath.scala 150:39:Sodor3Stage.fir@1347.4]
  assign _T_1005 = _T_1003 == 1'h0; // @[cpath.scala 150:25:Sodor3Stage.fir@1348.4]
  assign _T_1009 = io_imem_resp_valid == 1'h0; // @[cpath.scala 159:29:Sodor3Stage.fir@1359.4]
  assign rs1_addr = io_imem_resp_bits_inst[19:15]; // @[cpath.scala 162:41:Sodor3Stage.fir@1365.4]
  assign _T_1014 = cs0_7 == 3'h2; // @[cpath.scala 163:30:Sodor3Stage.fir@1366.4]
  assign _T_1015 = cs0_7 == 3'h3; // @[cpath.scala 163:54:Sodor3Stage.fir@1367.4]
  assign _T_1016 = _T_1014 | _T_1015; // @[cpath.scala 163:40:Sodor3Stage.fir@1368.4]
  assign _T_1018 = rs1_addr == 5'h0; // @[cpath.scala 163:77:Sodor3Stage.fir@1369.4]
  assign csr_ren = _T_1016 & _T_1018; // @[cpath.scala 163:65:Sodor3Stage.fir@1370.4]
  assign csr_cmd = csr_ren ? 3'h5 : cs0_7; // @[cpath.scala 164:21:Sodor3Stage.fir@1371.4]
  assign _T_1025 = cs_inst_val == 1'h0; // @[cpath.scala 178:24:Sodor3Stage.fir@1380.4]
  assign io_imem_req_valid = _T_1005 & io_imem_resp_valid;
  assign io_ctl_exe_kill = _T_1028 | io_dat_csr_eret;
  assign io_ctl_pc_sel = take_evec ? 3'h4 : _T_1002;
  assign io_ctl_brjmp_sel = _T_89 ? 1'h0 : _T_432;
  assign io_ctl_op1_sel = _T_89 ? 2'h0 : _T_481;
  assign io_ctl_op2_sel = _T_89 ? 2'h1 : _T_530;
  assign io_ctl_alu_fun = _T_89 ? 4'h0 : _T_579;
  assign io_ctl_wb_sel = _T_89 ? 2'h1 : _T_628;
  assign io_ctl_rf_wen = _T_1009 ? 1'h0 : cs0_2;
  assign io_ctl_bypassable = _T_89 ? 1'h0 : _T_726;
  assign io_ctl_csr_cmd = _T_1009 ? 3'h0 : csr_cmd;
  assign io_ctl_dmem_fcn = _T_89 ? 1'h0 : _T_824;
  assign io_ctl_dmem_typ = _T_89 ? 3'h3 : _T_873;
  assign io_ctl_exception = _T_1025 & io_imem_resp_valid;
  assign _GEN_91_0 = 32'h7033 == _T_164;
  assign _GEN_51_0 = 32'h7063 == _T_88;
  assign _GEN_304_0 = 32'h17 == _T_120;
  assign _GEN_199_0 = 32'h67 == _T_88;
  assign _GEN_148_0 = 32'h37 == _T_120;
  assign _GEN_403_0 = io_dat_br_eq;
  assign _GEN_24_0 = 32'h7033 == _T_164;
  assign _GEN_247_0 = 32'h7033 == _T_164;
  assign _GEN_106_0 = 32'h37 == _T_120;
  assign _GEN_133_0 = 32'h7033 == _T_164;
  assign _GEN_205_0 = 32'h7033 == _T_164;
  assign _GEN_39_0 = 32'h37 == _T_120;
  assign _GEN_232_0 = 32'h1073 == _T_88;
  assign _GEN_418_0 = _T_1016 & _T_1018;
  assign _GEN_127_0 = 32'h67 == _T_88;
  assign _GEN_331_0 = 32'h13 == _T_88;
  assign _GEN_190_0 = 32'h1073 == _T_88;
  assign _GEN_226_0 = 32'h1003 == _T_88;
  assign _GEN_45_0 = 32'h1003 == _T_88;
  assign _GEN_112_0 = 32'h1003 == _T_88;
  assign _GEN_298_0 = 32'h2013 == _T_88;
  assign _GEN_72_0 = 32'h4013 == _T_88;
  assign _GEN_211_0 = 32'h5013 == _T_152;
  assign _GEN_325_0 = 32'h1013 == _T_152;
  assign _GEN_397_0 = 32'h5003 == _T_88;
  assign _GEN_424_0 = 32'h2003 == _T_88;
  assign _GEN_30_0 = 32'h5013 == _T_152;
  assign _GEN_310_0 = 32'h4003 == _T_88;
  assign _GEN_319_0 = 32'h2033 == _T_164;
  assign _GEN_66_0 = 32'h1033 == _T_164;
  assign _GEN_220_0 = 32'h37 == _T_120;
  assign _GEN_214_0 = 32'h3013 == _T_88;
  assign _GEN_100_0 = 32'h3013 == _T_88;
  assign _GEN_109_0 = 32'h23 == _T_88;
  assign _GEN_313_0 = 32'h5033 == _T_164;
  assign _GEN_282_0 = 32'h67 == _T_88;
  assign _GEN_177_0 = 32'h13 == _T_88;
  assign _GEN_208_0 = 32'h40000033 == _T_164;
  assign _GEN_391_0 = 32'h13 == _T_88;
  assign _GEN_381_0 = 32'h33 == _T_164;
  assign _GEN_412_0 = cs_br_type == 4'h4;
  assign _GEN_27_0 = 32'h40000033 == _T_164;
  assign _GEN_276_0 = 32'h6063 == _T_88;
  assign _GEN_54_0 = 32'h63 == _T_88;
  assign _GEN_193_0 = 32'h6063 == _T_88;
  assign _GEN_12_1 = 32'h6063 == _T_88;
  assign _GEN_406_0 = io_dat_br_lt;
  assign _GEN_48_0 = 32'h2003 == _T_88;
  assign _GEN_115_0 = 32'h7073 == _T_88;
  assign _GEN_6_1 = 32'h7073 == _T_88;
  assign _GEN_33_0 = 32'h3013 == _T_88;
  assign _GEN_121_0 = 32'h6063 == _T_88;
  assign _GEN_307_0 = 32'h2023 == _T_88;
  assign _GEN_375_0 = 32'h4033 == _T_164;
  assign _GEN_229_0 = 32'h7073 == _T_88;
  assign _GEN_94_0 = 32'h40000033 == _T_164;
  assign _GEN_292_0 = 32'h33 == _T_164;
  assign _GEN_183_0 = 32'h5003 == _T_88;
  assign _GEN_0_1 = 32'h100f == _T_88;
  assign _GEN_196_0 = 32'h5063 == _T_88;
  assign _GEN_186_0 = 32'h3 == _T_88;
  assign _GEN_400_0 = 32'h3 == _T_88;
  assign _GEN_103_0 = 32'h6013 == _T_88;
  assign _GEN_264_0 = 32'h1023 == _T_88;
  assign _GEN_295_0 = 32'h40005013 == _T_152;
  assign _GEN_159_0 = 32'h5033 == _T_164;
  assign _GEN_202_0 = 32'h40005033 == _T_164;
  assign _GEN_171_0 = 32'h1013 == _T_152;
  assign _GEN_357_0 = 32'h30200073 == io_imem_resp_bits_inst;
  assign _GEN_270_0 = 32'h3 == _T_88;
  assign _GEN_384_0 = 32'h40005013 == _T_152;
  assign _GEN_36_0 = 32'h6013 == _T_88;
  assign _GEN_285_0 = 32'h40005033 == _T_164;
  assign _GEN_165_0 = 32'h2033 == _T_164;
  assign _GEN_279_0 = 32'h5063 == _T_88;
  assign _GEN_378_0 = 32'h3033 == _T_164;
  assign _GEN_21_1 = 32'h40005033 == _T_164;
  assign _GEN_301_0 = 32'h7013 == _T_88;
  assign _GEN_394_0 = 32'h1023 == _T_88;
  assign _GEN_15_1 = 32'h5063 == _T_88;
  assign _GEN_363_0 = 32'h6073 == _T_88;
  assign _GEN_9_3 = 32'h1073 == _T_88;
  assign _GEN_258_0 = 32'h4013 == _T_88;
  assign _GEN_97_0 = 32'h5013 == _T_152;
  assign _GEN_345_0 = 32'h4003 == _T_88;
  assign _GEN_339_0 = 32'h4003 == _T_88;
  assign _GEN_18_0 = 32'h67 == _T_88;
  assign _GEN_147_0 = 32'h13 == _T_88;
  assign _GEN_330_0 = 32'h7013 == _T_88;
  assign _GEN_86_0 = 32'h6f == _T_120;
  assign _GEN_273_0 = 32'h1073 == _T_88;
  assign _GEN_351_0 = 32'h1003 == _T_88;
  assign _GEN_231_0 = 32'h2073 == _T_88;
  assign _GEN_189_0 = 32'h2073 == _T_88;
  assign _GEN_153_0 = 32'h5003 == _T_88;
  assign _GEN_288_0 = 32'h7033 == _T_164;
  assign _GEN_366_0 = 32'h4063 == _T_88;
  assign _GEN_252_0 = 32'h1033 == _T_164;
  assign _GEN_180_0 = 32'h1023 == _T_88;
  assign _GEN_71_0 = 32'h2013 == _T_88;
  assign _GEN_174_0 = 32'h4013 == _T_88;
  assign _GEN_168_0 = 32'h1033 == _T_164;
  assign _GEN_372_0 = 32'h6f == _T_120;
  assign _GEN_3_2 = 32'h7b200073 == io_imem_resp_bits_inst;
  assign _GEN_387_0 = 32'h2013 == _T_88;
  assign _GEN_246_0 = 32'h6033 == _T_164;
  assign _GEN_267_0 = 32'h5003 == _T_88;
  assign _GEN_354_0 = 32'h10500073 == io_imem_resp_bits_inst;
  assign _GEN_213_0 = 32'h1013 == _T_152;
  assign _GEN_249_0 = 32'h2033 == _T_164;
  assign _GEN_240_0 = 32'h63 == _T_88;
  assign _GEN_141_0 = 32'h1013 == _T_152;
  assign _GEN_135_0 = 32'h2033 == _T_164;
  assign _GEN_234_0 = 32'h5073 == _T_88;
  assign _GEN_348_0 = 32'h23 == _T_88;
  assign _GEN_261_0 = 32'h13 == _T_88;
  assign _GEN_312_0 = 32'h2003 == _T_88;
  assign _GEN_53_0 = 32'h1063 == _T_88;
  assign _GEN_333_0 = 32'h17 == _T_120;
  assign _GEN_68_0 = 32'h40005013 == _T_152;
  assign _GEN_156_0 = 32'h3 == _T_88;
  assign _GEN_360_0 = 32'h3073 == _T_88;
  assign _GEN_369_0 = 32'h1063 == _T_88;
  assign _GEN_74_0 = 32'h7013 == _T_88;
  assign _GEN_327_0 = 32'h2013 == _T_88;
  assign _GEN_89_0 = 32'h4033 == _T_164;
  assign _GEN_162_0 = 32'h6033 == _T_164;
  assign _GEN_426_0 = 32'h2003 == _T_88;
  assign _GEN_129_0 = 32'h5033 == _T_164;
  assign _GEN_228_0 = 32'h3 == _T_88;
  assign _GEN_411_0 = cs_br_type == 4'h5;
  assign _GEN_255_0 = 32'h1013 == _T_152;
  assign _GEN_120_0 = 32'h5073 == _T_88;
  assign _GEN_80_0 = 32'h2023 == _T_88;
  assign _GEN_342_0 = 32'h2023 == _T_88;
  assign _GEN_393_0 = 32'h17 == _T_120;
  assign _GEN_56_0 = 32'h6f == _T_120;
  assign _GEN_144_0 = 32'h4013 == _T_88;
  assign _GEN_408_0 = cs_br_type == 4'h8;
  assign _GEN_222_0 = 32'h1023 == _T_88;
  assign _GEN_117_0 = 32'h2073 == _T_88;
  assign _GEN_321_0 = 32'h33 == _T_164;
  assign _GEN_243_0 = 32'h5033 == _T_164;
  assign _GEN_237_0 = 32'h7063 == _T_88;
  assign _GEN_123_0 = 32'h7063 == _T_88;
  assign _GEN_102_0 = 32'h4013 == _T_88;
  assign _GEN_62_0 = 32'h3033 == _T_164;
  assign _GEN_150_0 = 32'h1023 == _T_88;
  assign _GEN_336_0 = 32'h2023 == _T_88;
  assign _GEN_201_0 = 32'h5033 == _T_164;
  assign _GEN_195_0 = 32'h7063 == _T_88;
  assign _GEN_414_0 = cs_br_type == 4'h2;
  assign _GEN_300_0 = 32'h6013 == _T_88;
  assign _GEN_294_0 = 32'h5013 == _T_152;
  assign _GEN_309_0 = 32'h1003 == _T_88;
  assign _GEN_77_0 = 32'h17 == _T_120;
  assign _GEN_83_0 = 32'h4003 == _T_88;
  assign _GEN_216_0 = 32'h4013 == _T_88;
  assign _GEN_420_0 = 32'h2003 == _T_88;
  assign _GEN_35_0 = 32'h4013 == _T_88;
  assign _GEN_41_0 = 32'h1023 == _T_88;
  assign _GEN_315_0 = 32'h4033 == _T_164;
  assign _GEN_429_0 = 32'h2003 == _T_88;
  assign _GEN_138_0 = 32'h1033 == _T_164;
  assign _GEN_402_0 = io_dat_br_eq == 1'h0;
  assign _GEN_17_1 = 32'h63 == _T_88;
  assign _GEN_225_0 = 32'h5003 == _T_88;
  assign _GEN_105_0 = 32'h13 == _T_88;
  assign _GEN_50_0 = 32'h4063 == _T_88;
  assign _GEN_44_0 = 32'h5003 == _T_88;
  assign _GEN_324_0 = 32'h40005013 == _T_152;
  assign _GEN_318_0 = 32'h3033 == _T_164;
  assign _GEN_396_0 = 32'h2023 == _T_88;
  assign _GEN_386_0 = 32'h3013 == _T_88;
  assign _GEN_38_0 = 32'h13 == _T_88;
  assign _GEN_65_0 = 32'h33 == _T_164;
  assign _GEN_23_1 = 32'h6033 == _T_164;
  assign _GEN_417_0 = _T_1028 | io_dat_csr_eret;
  assign _GEN_111_0 = 32'h5003 == _T_88;
  assign _GEN_210_0 = 32'h1033 == _T_164;
  assign _GEN_219_0 = 32'h13 == _T_88;
  assign _GEN_423_0 = 32'h2003 == _T_88;
  assign _GEN_132_0 = 32'h6033 == _T_164;
  assign _GEN_126_0 = 32'h63 == _T_88;
  assign _GEN_287_0 = 32'h6033 == _T_164;
  assign _GEN_90_0 = 32'h6033 == _T_164;
  assign _GEN_204_0 = 32'h6033 == _T_164;
  assign _GEN_99_0 = 32'h1013 == _T_152;
  assign _GEN_303_0 = 32'h37 == _T_120;
  assign _GEN_297_0 = 32'h3013 == _T_88;
  assign _GEN_59_0 = 32'h4033 == _T_164;
  assign _GEN_188_0 = 32'h3073 == _T_88;
  assign _GEN_198_0 = 32'h63 == _T_88;
  assign _GEN_176_0 = 32'h7013 == _T_88;
  assign _GEN_11_3 = 32'h5073 == _T_88;
  assign _GEN_380_0 = 32'h40000033 == _T_164;
  assign _GEN_93_0 = 32'h2033 == _T_164;
  assign _GEN_161_0 = 32'h4033 == _T_164;
  assign _GEN_192_0 = 32'h5073 == _T_88;
  assign _GEN_207_0 = 32'h2033 == _T_164;
  assign _GEN_405_0 = io_dat_br_ltu == 1'h0;
  assign _GEN_260_0 = 32'h7013 == _T_88;
  assign _GEN_26_0 = 32'h2033 == _T_164;
  assign _GEN_114_0 = 32'h3 == _T_88;
  assign _GEN_269_0 = 32'h4003 == _T_88;
  assign _GEN_182_0 = 32'h2023 == _T_88;
  assign _GEN_399_0 = 32'h4003 == _T_88;
  assign _GEN_368_0 = 32'h5063 == _T_88;
  assign _GEN_390_0 = 32'h7013 == _T_88;
  assign _GEN_32_0 = 32'h1013 == _T_152;
  assign _GEN_281_0 = 32'h63 == _T_88;
  assign _GEN_275_0 = 32'h5073 == _T_88;
  assign _GEN_291_0 = 32'h40000033 == _T_164;
  assign _GEN_47_0 = 32'h3 == _T_88;
  assign _GEN_5_3 = 32'h73 == io_imem_resp_bits_inst;
  assign _GEN_389_0 = 32'h6013 == _T_88;
  assign _GEN_306_0 = 32'h23 == _T_88;
  assign _GEN_374_0 = 32'h40005033 == _T_164;
  assign _GEN_108_0 = 32'h1023 == _T_88;
  assign _GEN_356_0 = 32'h7b200073 == io_imem_resp_bits_inst;
  assign _GEN_20_1 = 32'h5033 == _T_164;
  assign _GEN_14_2 = 32'h7063 == _T_88;
  assign _GEN_29_0 = 32'h1033 == _T_164;
  assign _GEN_82_0 = 32'h1003 == _T_88;
  assign _GEN_170_0 = 32'h40005013 == _T_152;
  assign _GEN_185_0 = 32'h4003 == _T_88;
  assign _GEN_278_0 = 32'h7063 == _T_88;
  assign _GEN_143_0 = 32'h2013 == _T_88;
  assign _GEN_96_0 = 32'h1033 == _T_164;
  assign _GEN_263_0 = 32'h17 == _T_120;
  assign _GEN_164_0 = 32'h3033 == _T_164;
  assign _GEN_158_0 = 32'h6f == _T_120;
  assign _GEN_362_0 = 32'h1073 == _T_88;
  assign _GEN_377_0 = 32'h7033 == _T_164;
  assign _GEN_257_0 = 32'h2013 == _T_88;
  assign _GEN_284_0 = 32'h5033 == _T_164;
  assign _GEN_179_0 = 32'h17 == _T_120;
  assign _GEN_383_0 = 32'h5013 == _T_152;
  assign _GEN_242_0 = 32'h6f == _T_120;
  assign _GEN_8_3 = 32'h2073 == _T_88;
  assign _GEN_341_0 = 32'h23 == _T_88;
  assign _GEN_76_0 = 32'h37 == _T_120;
  assign _GEN_173_0 = 32'h2013 == _T_88;
  assign _GEN_224_1 = 32'h2023 == _T_88;
  assign _GEN_359_0 = 32'h7073 == _T_88;
  assign _GEN_251_0 = 32'h33 == _T_164;
  assign _GEN_131_0 = 32'h4033 == _T_164;
  assign _GEN_146_0 = 32'h7013 == _T_88;
  assign _GEN_350_0 = 32'h5003 == _T_88;
  assign _GEN_344_0 = 32'h1003 == _T_88;
  assign _GEN_239_1 = 32'h1063 == _T_88;
  assign _GEN_272_0 = 32'h2073 == _T_88;
  assign _GEN_64_0 = 32'h40000033 == _T_164;
  assign _GEN_58_0 = 32'h40005033 == _T_164;
  assign _GEN_230_0 = 32'h3073 == _T_88;
  assign _GEN_365_0 = 32'h6063 == _T_88;
  assign _GEN_323_1 = 32'h5013 == _T_152;
  assign _GEN_85_0 = 32'h2003 == _T_88;
  assign _GEN_338_1 = 32'h1003 == _T_88;
  assign _GEN_79_0 = 32'h23 == _T_88;
  assign _GEN_2_3 = 32'h100073 == io_imem_resp_bits_inst;
  assign _GEN_245_0 = 32'h4033 == _T_164;
  assign _GEN_70_0 = 32'h3013 == _T_88;
  assign _GEN_152_0 = 32'h2023 == _T_88;
  assign _GEN_167_0 = 32'h33 == _T_164;
  assign _GEN_422_0 = 32'h2003 == _T_88;
  assign _GEN_371_0 = 32'h67 == _T_88;
  assign _GEN_266_0 = 32'h2023 == _T_88;
  assign _GEN_125_0 = 32'h1063 == _T_88;
  assign _GEN_212_1 = 32'h40005013 == _T_152;
  assign _GEN_254_0 = 32'h40005013 == _T_152;
  assign _GEN_155_0 = 32'h4003 == _T_88;
  assign _GEN_149_0 = 32'h17 == _T_120;
  assign _GEN_227_0 = 32'h4003 == _T_88;
  assign _GEN_113_0 = 32'h4003 == _T_88;
  assign _GEN_140_0 = 32'h40005013 == _T_152;
  assign _GEN_326_0 = 32'h3013 == _T_88;
  assign _GEN_425_0 = io_imem_resp_valid == 1'h0;
  assign _GEN_404_0 = io_dat_br_lt == 1'h0;
  assign _GEN_353_0 = 32'h3 == _T_88;
  assign _GEN_248_0 = 32'h3033 == _T_164;
  assign _GEN_107_0 = 32'h17 == _T_120;
  assign _GEN_311_1 = 32'h3 == _T_88;
  assign _GEN_73_0 = 32'h6013 == _T_88;
  assign _GEN_67_0 = 32'h5013 == _T_152;
  assign _GEN_347_0 = 32'h1023 == _T_88;
  assign _GEN_206_1 = 32'h3033 == _T_164;
  assign _GEN_410_0 = cs_br_type == 4'h6;
  assign _GEN_419_0 = _T_1028 | io_dat_csr_eret;
  assign _GEN_233_0 = 32'h6073 == _T_88;
  assign _GEN_305_1 = 32'h1023 == _T_88;
  assign _GEN_128_0 = 32'h6f == _T_120;
  assign _GEN_332_0 = 32'h37 == _T_120;
  assign _GEN_88_0 = 32'h40005033 == _T_164;
  assign _GEN_52_0 = 32'h5063 == _T_88;
  assign _GEN_46_0 = 32'h4003 == _T_88;
  assign _GEN_134_0 = 32'h3033 == _T_164;
  assign _GEN_221_0 = 32'h17 == _T_120;
  assign _GEN_407_0 = io_dat_br_ltu;
  assign _GEN_382_1 = 32'h1033 == _T_164;
  assign _GEN_28_0 = 32'h33 == _T_164;
  assign _GEN_40_0 = 32'h17 == _T_120;
  assign _GEN_55_0 = 32'h67 == _T_88;
  assign _GEN_329_0 = 32'h6013 == _T_88;
  assign _GEN_194_1 = 32'h4063 == _T_88;
  assign _GEN_392_0 = 32'h37 == _T_120;
  assign _GEN_236_0 = 32'h4063 == _T_88;
  assign _GEN_101_0 = 32'h2013 == _T_88;
  assign _GEN_61_0 = 32'h7033 == _T_164;
  assign _GEN_34_0 = 32'h2013 == _T_88;
  assign _GEN_116_0 = 32'h3073 == _T_88;
  assign _GEN_122_0 = 32'h4063 == _T_88;
  assign _GEN_320_1 = 32'h40000033 == _T_164;
  assign _GEN_215_0 = 32'h2013 == _T_88;
  assign _GEN_335_0 = 32'h23 == _T_88;
  assign _GEN_293_1 = 32'h1033 == _T_164;
  assign _GEN_428_0 = 32'h2003 == _T_88;
  assign _GEN_49_0 = 32'h6063 == _T_88;
  assign _GEN_137_0 = 32'h33 == _T_164;
  assign _GEN_200_1 = 32'h6f == _T_120;
  assign _GEN_209_0 = 32'h33 == _T_164;
  assign _GEN_95_0 = 32'h33 == _T_164;
  assign _GEN_413_0 = cs_br_type == 4'h3;
  assign _GEN_314_0 = 32'h40005033 == _T_164;
  assign _GEN_308_0 = 32'h5003 == _T_88;
  assign _GEN_16_1 = 32'h1063 == _T_88;
  assign _GEN_395_0 = 32'h23 == _T_88;
  assign _GEN_385_1 = 32'h1013 == _T_152;
  assign _GEN_104_0 = 32'h7013 == _T_88;
  assign _GEN_302_1 = 32'h13 == _T_88;
  assign _GEN_317_1 = 32'h7033 == _T_164;
  assign _GEN_203_1 = 32'h4033 == _T_164;
  assign _GEN_172_1 = 32'h3013 == _T_88;
  assign _GEN_197_1 = 32'h1063 == _T_88;
  assign _GEN_370_1 = 32'h63 == _T_88;
  assign _GEN_416_0 = cs_br_type == 4'h0;
  assign _GEN_22_1 = 32'h4033 == _T_164;
  assign _GEN_271_1 = 32'h3073 == _T_88;
  assign _GEN_119_0 = 32'h6073 == _T_88;
  assign _GEN_379_1 = 32'h2033 == _T_164;
  assign _GEN_187_1 = 32'h7073 == _T_88;
  assign _GEN_401_0 = 32'h2003 == _T_88;
  assign _GEN_43_0 = 32'h2023 == _T_88;
  assign _GEN_296_1 = 32'h1013 == _T_152;
  assign _GEN_286_1 = 32'h4033 == _T_164;
  assign _GEN_364_1 = 32'h5073 == _T_88;
  assign _GEN_1_5 = 32'h10500073 == io_imem_resp_bits_inst;
  assign _GEN_98_0 = 32'h40005013 == _T_152;
  assign _GEN_37_0 = 32'h7013 == _T_88;
  assign _GEN_110_0 = 32'h2023 == _T_88;
  assign _GEN_218_1 = 32'h7013 == _T_88;
  assign _GEN_25_0 = 32'h3033 == _T_164;
  assign _GEN_181_1 = 32'h23 == _T_88;
  assign _GEN_175_1 = 32'h6013 == _T_88;
  assign _GEN_289_1 = 32'h3033 == _T_164;
  assign _GEN_352_1 = 32'h4003 == _T_88;
  assign _GEN_31_0 = 32'h40005013 == _T_152;
  assign _GEN_274_1 = 32'h6073 == _T_88;
  assign _GEN_160_1 = 32'h40005033 == _T_164;
  assign _GEN_169_1 = 32'h5013 == _T_152;
  assign _GEN_191_1 = 32'h6073 == _T_88;
  assign _GEN_373_1 = 32'h5033 == _T_164;
  assign _GEN_19_1 = 32'h6f == _T_120;
  assign _GEN_367_1 = 32'h7063 == _T_88;
  assign _GEN_268_1 = 32'h1003 == _T_88;
  assign _GEN_290_1 = 32'h2033 == _T_164;
  assign _GEN_280_1 = 32'h1063 == _T_88;
  assign _GEN_154_1 = 32'h1003 == _T_88;
  assign _GEN_87_0 = 32'h5033 == _T_164;
  assign _GEN_299_1 = 32'h4013 == _T_88;
  assign _GEN_10_4 = 32'h6073 == _T_88;
  assign _GEN_398_0 = 32'h1003 == _T_88;
  assign _GEN_4_4 = 32'h30200073 == io_imem_resp_bits_inst;
  assign _GEN_388_1 = 32'h4013 == _T_88;
  assign _GEN_253_1 = 32'h5013 == _T_152;
  assign _GEN_92_0 = 32'h3033 == _T_164;
  assign _GEN_346_1 = 32'h3 == _T_88;
  assign _GEN_334_1 = 32'h1023 == _T_88;
  assign _GEN_340_1 = 32'h3 == _T_88;
  assign _GEN_13_3 = 32'h4063 == _T_88;
  assign _GEN_256_1 = 32'h3013 == _T_88;
  assign _GEN_328_1 = 32'h4013 == _T_88;
  assign _GEN_81_0 = 32'h5003 == _T_88;
  assign _GEN_355_1 = 32'h100073 == io_imem_resp_bits_inst;
  assign _GEN_7_6 = 32'h3073 == _T_88;
  assign _GEN_277_1 = 32'h4063 == _T_88;
  assign _GEN_69_0 = 32'h1013 == _T_152;
  assign _GEN_157_1 = 32'h67 == _T_88;
  assign _GEN_235_1 = 32'h6063 == _T_88;
  assign _GEN_184_1 = 32'h1003 == _T_88;
  assign _GEN_60_0 = 32'h6033 == _T_164;
  assign _GEN_283_1 = 32'h6f == _T_120;
  assign _GEN_142_0 = 32'h3013 == _T_88;
  assign _GEN_178_1 = 32'h37 == _T_120;
  assign _GEN_241_1 = 32'h67 == _T_88;
  assign _GEN_361_1 = 32'h2073 == _T_88;
  assign _GEN_136_0 = 32'h40000033 == _T_164;
  assign _GEN_75_0 = 32'h13 == _T_88;
  assign _GEN_163_1 = 32'h7033 == _T_164;
  assign _GEN_349_1 = 32'h2023 == _T_88;
  assign _GEN_427_0 = io_imem_resp_valid == 1'h0;
  assign _GEN_376_1 = 32'h6033 == _T_164;
  assign _GEN_262_1 = 32'h37 == _T_120;
  assign _GEN_166_1 = 32'h40000033 == _T_164;
  assign _GEN_358_1 = 32'h73 == io_imem_resp_bits_inst;
  assign _GEN_42_0 = 32'h23 == _T_88;
  assign _GEN_265_1 = 32'h23 == _T_88;
  assign _GEN_316_1 = 32'h6033 == _T_164;
  assign _GEN_130_0 = 32'h40005033 == _T_164;
  assign _GEN_124_0 = 32'h5063 == _T_88;
  assign _GEN_343_1 = 32'h5003 == _T_88;
  assign _GEN_223_1 = 32'h23 == _T_88;
  assign _GEN_238_1 = 32'h5063 == _T_88;
  assign _GEN_118_0 = 32'h1073 == _T_88;
  assign _GEN_151_1 = 32'h23 == _T_88;
  assign _GEN_145_0 = 32'h6013 == _T_88;
  assign _GEN_337_1 = 32'h5003 == _T_88;
  assign _GEN_244_1 = 32'h40005033 == _T_164;
  assign _GEN_409_0 = cs_br_type == 4'h7;
  assign _GEN_322_1 = 32'h1033 == _T_164;
  assign _GEN_78_0 = 32'h1023 == _T_88;
  assign _GEN_217_1 = 32'h6013 == _T_88;
  assign _GEN_421_0 = 32'h2003 == _T_88;
  assign _GEN_415_0 = cs_br_type == 4'h1;
  assign _GEN_63_0 = 32'h2033 == _T_164;
  assign _GEN_57_0 = 32'h5033 == _T_164;
  assign _GEN_250_1 = 32'h40000033 == _T_164;
  assign _GEN_259_1 = 32'h6013 == _T_88;
  assign _GEN_139_0 = 32'h5013 == _T_152;
  assign _GEN_84_0 = 32'h3 == _T_88;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_1028 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (metaReset) begin
      _T_1028 <= 1'h0;
    end else begin
      _T_1028 <= io_ctl_exception;
    end
  end
endmodule
module ALU( // @[:Sodor3Stage.fir@1388.2]
  input  [3:0]  io_fn, // @[:Sodor3Stage.fir@1391.4]
  input  [31:0] io_in2, // @[:Sodor3Stage.fir@1391.4]
  input  [31:0] io_in1, // @[:Sodor3Stage.fir@1391.4]
  output [31:0] io_out, // @[:Sodor3Stage.fir@1391.4]
  output [31:0] io_adder_out, // @[:Sodor3Stage.fir@1391.4]
  output        _GEN_9_1,
  output        _GEN_0_0,
  output        _GEN_8_0,
  output        _GEN_2_0,
  output        _GEN_5_1,
  output        _GEN_10_1,
  output        _GEN_7_2,
  output        _GEN_1_4,
  output        _GEN_4_2,
  output        _GEN_3_5,
  output        _GEN_6_5
);
  wire  _T_9; // @[alu.scala 30:29:Sodor3Stage.fir@1393.4]
  wire [32:0] _T_11; // @[alu.scala 50:40:Sodor3Stage.fir@1394.4]
  wire [32:0] _T_12; // @[alu.scala 50:40:Sodor3Stage.fir@1395.4]
  wire [31:0] _T_13; // @[alu.scala 50:40:Sodor3Stage.fir@1396.4]
  wire [31:0] _T_14; // @[alu.scala 50:25:Sodor3Stage.fir@1397.4]
  wire [32:0] _T_15; // @[alu.scala 50:20:Sodor3Stage.fir@1398.4]
  wire [31:0] sum; // @[alu.scala 50:20:Sodor3Stage.fir@1399.4]
  wire  _T_16; // @[alu.scala 53:26:Sodor3Stage.fir@1400.4]
  wire  _T_17; // @[alu.scala 53:42:Sodor3Stage.fir@1401.4]
  wire  _T_18; // @[alu.scala 53:32:Sodor3Stage.fir@1402.4]
  wire  _T_19; // @[alu.scala 53:52:Sodor3Stage.fir@1403.4]
  wire  _T_20; // @[alu.scala 31:30:Sodor3Stage.fir@1404.4]
  wire  _T_23; // @[alu.scala 54:18:Sodor3Stage.fir@1407.4]
  wire  less; // @[alu.scala 53:19:Sodor3Stage.fir@1408.4]
  wire [4:0] shamt; // @[alu.scala 58:21:Sodor3Stage.fir@1409.4]
  wire  _T_24; // @[alu.scala 60:24:Sodor3Stage.fir@1411.4]
  wire  _T_25; // @[alu.scala 60:46:Sodor3Stage.fir@1412.4]
  wire  _T_26; // @[alu.scala 60:37:Sodor3Stage.fir@1413.4]
  wire [15:0] _T_31; // @[Bitwise.scala 103:21:Sodor3Stage.fir@1416.4]
  wire [31:0] _T_32; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1417.4]
  wire [15:0] _T_33; // @[Bitwise.scala 103:46:Sodor3Stage.fir@1418.4]
  wire [31:0] _GEN_11; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1419.4]
  wire [31:0] _T_34; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1419.4]
  wire [31:0] _T_36; // @[Bitwise.scala 103:75:Sodor3Stage.fir@1421.4]
  wire [31:0] _T_37; // @[Bitwise.scala 103:39:Sodor3Stage.fir@1422.4]
  wire [23:0] _T_41; // @[Bitwise.scala 103:21:Sodor3Stage.fir@1426.4]
  wire [31:0] _GEN_12; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1427.4]
  wire [31:0] _T_42; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1427.4]
  wire [23:0] _T_43; // @[Bitwise.scala 103:46:Sodor3Stage.fir@1428.4]
  wire [31:0] _GEN_13; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1429.4]
  wire [31:0] _T_44; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1429.4]
  wire [31:0] _T_46; // @[Bitwise.scala 103:75:Sodor3Stage.fir@1431.4]
  wire [31:0] _T_47; // @[Bitwise.scala 103:39:Sodor3Stage.fir@1432.4]
  wire [27:0] _T_51; // @[Bitwise.scala 103:21:Sodor3Stage.fir@1436.4]
  wire [31:0] _GEN_14; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1437.4]
  wire [31:0] _T_52; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1437.4]
  wire [27:0] _T_53; // @[Bitwise.scala 103:46:Sodor3Stage.fir@1438.4]
  wire [31:0] _GEN_15; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1439.4]
  wire [31:0] _T_54; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1439.4]
  wire [31:0] _T_56; // @[Bitwise.scala 103:75:Sodor3Stage.fir@1441.4]
  wire [31:0] _T_57; // @[Bitwise.scala 103:39:Sodor3Stage.fir@1442.4]
  wire [29:0] _T_61; // @[Bitwise.scala 103:21:Sodor3Stage.fir@1446.4]
  wire [31:0] _GEN_16; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1447.4]
  wire [31:0] _T_62; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1447.4]
  wire [29:0] _T_63; // @[Bitwise.scala 103:46:Sodor3Stage.fir@1448.4]
  wire [31:0] _GEN_17; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1449.4]
  wire [31:0] _T_64; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1449.4]
  wire [31:0] _T_66; // @[Bitwise.scala 103:75:Sodor3Stage.fir@1451.4]
  wire [31:0] _T_67; // @[Bitwise.scala 103:39:Sodor3Stage.fir@1452.4]
  wire [30:0] _T_71; // @[Bitwise.scala 103:21:Sodor3Stage.fir@1456.4]
  wire [31:0] _GEN_18; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1457.4]
  wire [31:0] _T_72; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1457.4]
  wire [30:0] _T_73; // @[Bitwise.scala 103:46:Sodor3Stage.fir@1458.4]
  wire [31:0] _GEN_19; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1459.4]
  wire [31:0] _T_74; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1459.4]
  wire [31:0] _T_76; // @[Bitwise.scala 103:75:Sodor3Stage.fir@1461.4]
  wire [31:0] _T_77; // @[Bitwise.scala 103:39:Sodor3Stage.fir@1462.4]
  wire [31:0] shin; // @[alu.scala 60:17:Sodor3Stage.fir@1463.4]
  wire  _T_79; // @[alu.scala 61:41:Sodor3Stage.fir@1465.4]
  wire  _T_80; // @[alu.scala 61:35:Sodor3Stage.fir@1466.4]
  wire [32:0] _T_81; // @[Cat.scala 30:58:Sodor3Stage.fir@1467.4]
  wire [32:0] _T_82; // @[:Sodor3Stage.fir@1468.4]
  wire [32:0] _T_83; // @[alu.scala 61:61:Sodor3Stage.fir@1469.4]
  wire [31:0] shout_r; // @[alu.scala 61:70:Sodor3Stage.fir@1470.4]
  wire [15:0] _T_88; // @[Bitwise.scala 103:21:Sodor3Stage.fir@1473.4]
  wire [31:0] _T_89; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1474.4]
  wire [15:0] _T_90; // @[Bitwise.scala 103:46:Sodor3Stage.fir@1475.4]
  wire [31:0] _GEN_20; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1476.4]
  wire [31:0] _T_91; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1476.4]
  wire [31:0] _T_93; // @[Bitwise.scala 103:75:Sodor3Stage.fir@1478.4]
  wire [31:0] _T_94; // @[Bitwise.scala 103:39:Sodor3Stage.fir@1479.4]
  wire [23:0] _T_98; // @[Bitwise.scala 103:21:Sodor3Stage.fir@1483.4]
  wire [31:0] _GEN_21; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1484.4]
  wire [31:0] _T_99; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1484.4]
  wire [23:0] _T_100; // @[Bitwise.scala 103:46:Sodor3Stage.fir@1485.4]
  wire [31:0] _GEN_22; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1486.4]
  wire [31:0] _T_101; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1486.4]
  wire [31:0] _T_103; // @[Bitwise.scala 103:75:Sodor3Stage.fir@1488.4]
  wire [31:0] _T_104; // @[Bitwise.scala 103:39:Sodor3Stage.fir@1489.4]
  wire [27:0] _T_108; // @[Bitwise.scala 103:21:Sodor3Stage.fir@1493.4]
  wire [31:0] _GEN_23; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1494.4]
  wire [31:0] _T_109; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1494.4]
  wire [27:0] _T_110; // @[Bitwise.scala 103:46:Sodor3Stage.fir@1495.4]
  wire [31:0] _GEN_24; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1496.4]
  wire [31:0] _T_111; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1496.4]
  wire [31:0] _T_113; // @[Bitwise.scala 103:75:Sodor3Stage.fir@1498.4]
  wire [31:0] _T_114; // @[Bitwise.scala 103:39:Sodor3Stage.fir@1499.4]
  wire [29:0] _T_118; // @[Bitwise.scala 103:21:Sodor3Stage.fir@1503.4]
  wire [31:0] _GEN_25; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1504.4]
  wire [31:0] _T_119; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1504.4]
  wire [29:0] _T_120; // @[Bitwise.scala 103:46:Sodor3Stage.fir@1505.4]
  wire [31:0] _GEN_26; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1506.4]
  wire [31:0] _T_121; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1506.4]
  wire [31:0] _T_123; // @[Bitwise.scala 103:75:Sodor3Stage.fir@1508.4]
  wire [31:0] _T_124; // @[Bitwise.scala 103:39:Sodor3Stage.fir@1509.4]
  wire [30:0] _T_128; // @[Bitwise.scala 103:21:Sodor3Stage.fir@1513.4]
  wire [31:0] _GEN_27; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1514.4]
  wire [31:0] _T_129; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1514.4]
  wire [30:0] _T_130; // @[Bitwise.scala 103:46:Sodor3Stage.fir@1515.4]
  wire [31:0] _GEN_28; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1516.4]
  wire [31:0] _T_131; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1516.4]
  wire [31:0] _T_133; // @[Bitwise.scala 103:75:Sodor3Stage.fir@1518.4]
  wire [31:0] shout_l; // @[Bitwise.scala 103:39:Sodor3Stage.fir@1519.4]
  wire  _T_134; // @[alu.scala 65:15:Sodor3Stage.fir@1520.4]
  wire [31:0] _T_135; // @[alu.scala 65:35:Sodor3Stage.fir@1521.4]
  wire  _T_136; // @[alu.scala 66:15:Sodor3Stage.fir@1522.4]
  wire [31:0] _T_137; // @[alu.scala 66:35:Sodor3Stage.fir@1523.4]
  wire  _T_138; // @[alu.scala 67:15:Sodor3Stage.fir@1524.4]
  wire [31:0] _T_139; // @[alu.scala 67:35:Sodor3Stage.fir@1525.4]
  wire [31:0] _T_140; // @[alu.scala 67:8:Sodor3Stage.fir@1526.4]
  wire [31:0] _T_141; // @[alu.scala 66:8:Sodor3Stage.fir@1527.4]
  wire [31:0] bitwise_logic; // @[alu.scala 65:8:Sodor3Stage.fir@1528.4]
  wire  _T_142; // @[alu.scala 71:15:Sodor3Stage.fir@1529.4]
  wire  _T_143; // @[alu.scala 71:36:Sodor3Stage.fir@1530.4]
  wire  _T_144; // @[alu.scala 71:27:Sodor3Stage.fir@1531.4]
  wire  _T_145; // @[alu.scala 72:15:Sodor3Stage.fir@1532.4]
  wire  _T_146; // @[alu.scala 72:36:Sodor3Stage.fir@1533.4]
  wire  _T_147; // @[alu.scala 72:27:Sodor3Stage.fir@1534.4]
  wire  _T_151; // @[alu.scala 74:15:Sodor3Stage.fir@1538.4]
  wire [31:0] _T_152; // @[alu.scala 74:8:Sodor3Stage.fir@1539.4]
  wire [31:0] _T_153; // @[alu.scala 73:8:Sodor3Stage.fir@1540.4]
  wire [31:0] _T_154; // @[alu.scala 72:8:Sodor3Stage.fir@1541.4]
  assign _T_9 = io_fn[3]; // @[alu.scala 30:29:Sodor3Stage.fir@1393.4]
  assign _T_11 = 32'h0 - io_in2; // @[alu.scala 50:40:Sodor3Stage.fir@1394.4]
  assign _T_12 = $unsigned(_T_11); // @[alu.scala 50:40:Sodor3Stage.fir@1395.4]
  assign _T_13 = _T_12[31:0]; // @[alu.scala 50:40:Sodor3Stage.fir@1396.4]
  assign _T_14 = _T_9 ? _T_13 : io_in2; // @[alu.scala 50:25:Sodor3Stage.fir@1397.4]
  assign _T_15 = io_in1 + _T_14; // @[alu.scala 50:20:Sodor3Stage.fir@1398.4]
  assign sum = _T_15[31:0]; // @[alu.scala 50:20:Sodor3Stage.fir@1399.4]
  assign _T_16 = io_in1[31]; // @[alu.scala 53:26:Sodor3Stage.fir@1400.4]
  assign _T_17 = io_in2[31]; // @[alu.scala 53:42:Sodor3Stage.fir@1401.4]
  assign _T_18 = _T_16 == _T_17; // @[alu.scala 53:32:Sodor3Stage.fir@1402.4]
  assign _T_19 = sum[31]; // @[alu.scala 53:52:Sodor3Stage.fir@1403.4]
  assign _T_20 = io_fn[1]; // @[alu.scala 31:30:Sodor3Stage.fir@1404.4]
  assign _T_23 = _T_20 ? _T_17 : _T_16; // @[alu.scala 54:18:Sodor3Stage.fir@1407.4]
  assign less = _T_18 ? _T_19 : _T_23; // @[alu.scala 53:19:Sodor3Stage.fir@1408.4]
  assign shamt = io_in2[4:0]; // @[alu.scala 58:21:Sodor3Stage.fir@1409.4]
  assign _T_24 = io_fn == 4'h5; // @[alu.scala 60:24:Sodor3Stage.fir@1411.4]
  assign _T_25 = io_fn == 4'hb; // @[alu.scala 60:46:Sodor3Stage.fir@1412.4]
  assign _T_26 = _T_24 | _T_25; // @[alu.scala 60:37:Sodor3Stage.fir@1413.4]
  assign _T_31 = io_in1[31:16]; // @[Bitwise.scala 103:21:Sodor3Stage.fir@1416.4]
  assign _T_32 = {{16'd0}, _T_31}; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1417.4]
  assign _T_33 = io_in1[15:0]; // @[Bitwise.scala 103:46:Sodor3Stage.fir@1418.4]
  assign _GEN_11 = {{16'd0}, _T_33}; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1419.4]
  assign _T_34 = _GEN_11 << 16; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1419.4]
  assign _T_36 = _T_34 & 32'hffff0000; // @[Bitwise.scala 103:75:Sodor3Stage.fir@1421.4]
  assign _T_37 = _T_32 | _T_36; // @[Bitwise.scala 103:39:Sodor3Stage.fir@1422.4]
  assign _T_41 = _T_37[31:8]; // @[Bitwise.scala 103:21:Sodor3Stage.fir@1426.4]
  assign _GEN_12 = {{8'd0}, _T_41}; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1427.4]
  assign _T_42 = _GEN_12 & 32'hff00ff; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1427.4]
  assign _T_43 = _T_37[23:0]; // @[Bitwise.scala 103:46:Sodor3Stage.fir@1428.4]
  assign _GEN_13 = {{8'd0}, _T_43}; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1429.4]
  assign _T_44 = _GEN_13 << 8; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1429.4]
  assign _T_46 = _T_44 & 32'hff00ff00; // @[Bitwise.scala 103:75:Sodor3Stage.fir@1431.4]
  assign _T_47 = _T_42 | _T_46; // @[Bitwise.scala 103:39:Sodor3Stage.fir@1432.4]
  assign _T_51 = _T_47[31:4]; // @[Bitwise.scala 103:21:Sodor3Stage.fir@1436.4]
  assign _GEN_14 = {{4'd0}, _T_51}; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1437.4]
  assign _T_52 = _GEN_14 & 32'hf0f0f0f; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1437.4]
  assign _T_53 = _T_47[27:0]; // @[Bitwise.scala 103:46:Sodor3Stage.fir@1438.4]
  assign _GEN_15 = {{4'd0}, _T_53}; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1439.4]
  assign _T_54 = _GEN_15 << 4; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1439.4]
  assign _T_56 = _T_54 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75:Sodor3Stage.fir@1441.4]
  assign _T_57 = _T_52 | _T_56; // @[Bitwise.scala 103:39:Sodor3Stage.fir@1442.4]
  assign _T_61 = _T_57[31:2]; // @[Bitwise.scala 103:21:Sodor3Stage.fir@1446.4]
  assign _GEN_16 = {{2'd0}, _T_61}; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1447.4]
  assign _T_62 = _GEN_16 & 32'h33333333; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1447.4]
  assign _T_63 = _T_57[29:0]; // @[Bitwise.scala 103:46:Sodor3Stage.fir@1448.4]
  assign _GEN_17 = {{2'd0}, _T_63}; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1449.4]
  assign _T_64 = _GEN_17 << 2; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1449.4]
  assign _T_66 = _T_64 & 32'hcccccccc; // @[Bitwise.scala 103:75:Sodor3Stage.fir@1451.4]
  assign _T_67 = _T_62 | _T_66; // @[Bitwise.scala 103:39:Sodor3Stage.fir@1452.4]
  assign _T_71 = _T_67[31:1]; // @[Bitwise.scala 103:21:Sodor3Stage.fir@1456.4]
  assign _GEN_18 = {{1'd0}, _T_71}; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1457.4]
  assign _T_72 = _GEN_18 & 32'h55555555; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1457.4]
  assign _T_73 = _T_67[30:0]; // @[Bitwise.scala 103:46:Sodor3Stage.fir@1458.4]
  assign _GEN_19 = {{1'd0}, _T_73}; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1459.4]
  assign _T_74 = _GEN_19 << 1; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1459.4]
  assign _T_76 = _T_74 & 32'haaaaaaaa; // @[Bitwise.scala 103:75:Sodor3Stage.fir@1461.4]
  assign _T_77 = _T_72 | _T_76; // @[Bitwise.scala 103:39:Sodor3Stage.fir@1462.4]
  assign shin = _T_26 ? io_in1 : _T_77; // @[alu.scala 60:17:Sodor3Stage.fir@1463.4]
  assign _T_79 = shin[31]; // @[alu.scala 61:41:Sodor3Stage.fir@1465.4]
  assign _T_80 = _T_9 & _T_79; // @[alu.scala 61:35:Sodor3Stage.fir@1466.4]
  assign _T_81 = {_T_80,shin}; // @[Cat.scala 30:58:Sodor3Stage.fir@1467.4]
  assign _T_82 = $signed(_T_81); // @[:Sodor3Stage.fir@1468.4]
  assign _T_83 = $signed(_T_82) >>> shamt; // @[alu.scala 61:61:Sodor3Stage.fir@1469.4]
  assign shout_r = _T_83[31:0]; // @[alu.scala 61:70:Sodor3Stage.fir@1470.4]
  assign _T_88 = shout_r[31:16]; // @[Bitwise.scala 103:21:Sodor3Stage.fir@1473.4]
  assign _T_89 = {{16'd0}, _T_88}; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1474.4]
  assign _T_90 = shout_r[15:0]; // @[Bitwise.scala 103:46:Sodor3Stage.fir@1475.4]
  assign _GEN_20 = {{16'd0}, _T_90}; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1476.4]
  assign _T_91 = _GEN_20 << 16; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1476.4]
  assign _T_93 = _T_91 & 32'hffff0000; // @[Bitwise.scala 103:75:Sodor3Stage.fir@1478.4]
  assign _T_94 = _T_89 | _T_93; // @[Bitwise.scala 103:39:Sodor3Stage.fir@1479.4]
  assign _T_98 = _T_94[31:8]; // @[Bitwise.scala 103:21:Sodor3Stage.fir@1483.4]
  assign _GEN_21 = {{8'd0}, _T_98}; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1484.4]
  assign _T_99 = _GEN_21 & 32'hff00ff; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1484.4]
  assign _T_100 = _T_94[23:0]; // @[Bitwise.scala 103:46:Sodor3Stage.fir@1485.4]
  assign _GEN_22 = {{8'd0}, _T_100}; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1486.4]
  assign _T_101 = _GEN_22 << 8; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1486.4]
  assign _T_103 = _T_101 & 32'hff00ff00; // @[Bitwise.scala 103:75:Sodor3Stage.fir@1488.4]
  assign _T_104 = _T_99 | _T_103; // @[Bitwise.scala 103:39:Sodor3Stage.fir@1489.4]
  assign _T_108 = _T_104[31:4]; // @[Bitwise.scala 103:21:Sodor3Stage.fir@1493.4]
  assign _GEN_23 = {{4'd0}, _T_108}; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1494.4]
  assign _T_109 = _GEN_23 & 32'hf0f0f0f; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1494.4]
  assign _T_110 = _T_104[27:0]; // @[Bitwise.scala 103:46:Sodor3Stage.fir@1495.4]
  assign _GEN_24 = {{4'd0}, _T_110}; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1496.4]
  assign _T_111 = _GEN_24 << 4; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1496.4]
  assign _T_113 = _T_111 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75:Sodor3Stage.fir@1498.4]
  assign _T_114 = _T_109 | _T_113; // @[Bitwise.scala 103:39:Sodor3Stage.fir@1499.4]
  assign _T_118 = _T_114[31:2]; // @[Bitwise.scala 103:21:Sodor3Stage.fir@1503.4]
  assign _GEN_25 = {{2'd0}, _T_118}; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1504.4]
  assign _T_119 = _GEN_25 & 32'h33333333; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1504.4]
  assign _T_120 = _T_114[29:0]; // @[Bitwise.scala 103:46:Sodor3Stage.fir@1505.4]
  assign _GEN_26 = {{2'd0}, _T_120}; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1506.4]
  assign _T_121 = _GEN_26 << 2; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1506.4]
  assign _T_123 = _T_121 & 32'hcccccccc; // @[Bitwise.scala 103:75:Sodor3Stage.fir@1508.4]
  assign _T_124 = _T_119 | _T_123; // @[Bitwise.scala 103:39:Sodor3Stage.fir@1509.4]
  assign _T_128 = _T_124[31:1]; // @[Bitwise.scala 103:21:Sodor3Stage.fir@1513.4]
  assign _GEN_27 = {{1'd0}, _T_128}; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1514.4]
  assign _T_129 = _GEN_27 & 32'h55555555; // @[Bitwise.scala 103:31:Sodor3Stage.fir@1514.4]
  assign _T_130 = _T_124[30:0]; // @[Bitwise.scala 103:46:Sodor3Stage.fir@1515.4]
  assign _GEN_28 = {{1'd0}, _T_130}; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1516.4]
  assign _T_131 = _GEN_28 << 1; // @[Bitwise.scala 103:65:Sodor3Stage.fir@1516.4]
  assign _T_133 = _T_131 & 32'haaaaaaaa; // @[Bitwise.scala 103:75:Sodor3Stage.fir@1518.4]
  assign shout_l = _T_129 | _T_133; // @[Bitwise.scala 103:39:Sodor3Stage.fir@1519.4]
  assign _T_134 = io_fn == 4'h7; // @[alu.scala 65:15:Sodor3Stage.fir@1520.4]
  assign _T_135 = io_in1 & io_in2; // @[alu.scala 65:35:Sodor3Stage.fir@1521.4]
  assign _T_136 = io_fn == 4'h6; // @[alu.scala 66:15:Sodor3Stage.fir@1522.4]
  assign _T_137 = io_in1 | io_in2; // @[alu.scala 66:35:Sodor3Stage.fir@1523.4]
  assign _T_138 = io_fn == 4'h4; // @[alu.scala 67:15:Sodor3Stage.fir@1524.4]
  assign _T_139 = io_in1 ^ io_in2; // @[alu.scala 67:35:Sodor3Stage.fir@1525.4]
  assign _T_140 = _T_138 ? _T_139 : io_in1; // @[alu.scala 67:8:Sodor3Stage.fir@1526.4]
  assign _T_141 = _T_136 ? _T_137 : _T_140; // @[alu.scala 66:8:Sodor3Stage.fir@1527.4]
  assign bitwise_logic = _T_134 ? _T_135 : _T_141; // @[alu.scala 65:8:Sodor3Stage.fir@1528.4]
  assign _T_142 = io_fn == 4'h0; // @[alu.scala 71:15:Sodor3Stage.fir@1529.4]
  assign _T_143 = io_fn == 4'ha; // @[alu.scala 71:36:Sodor3Stage.fir@1530.4]
  assign _T_144 = _T_142 | _T_143; // @[alu.scala 71:27:Sodor3Stage.fir@1531.4]
  assign _T_145 = io_fn == 4'hc; // @[alu.scala 72:15:Sodor3Stage.fir@1532.4]
  assign _T_146 = io_fn == 4'he; // @[alu.scala 72:36:Sodor3Stage.fir@1533.4]
  assign _T_147 = _T_145 | _T_146; // @[alu.scala 72:27:Sodor3Stage.fir@1534.4]
  assign _T_151 = io_fn == 4'h1; // @[alu.scala 74:15:Sodor3Stage.fir@1538.4]
  assign _T_152 = _T_151 ? shout_l : bitwise_logic; // @[alu.scala 74:8:Sodor3Stage.fir@1539.4]
  assign _T_153 = _T_26 ? shout_r : _T_152; // @[alu.scala 73:8:Sodor3Stage.fir@1540.4]
  assign _T_154 = _T_147 ? {{31'd0}, less} : _T_153; // @[alu.scala 72:8:Sodor3Stage.fir@1541.4]
  assign io_out = _T_144 ? sum : _T_154;
  assign io_adder_out = _T_15[31:0];
  assign _GEN_9_1 = _T_145 | _T_146;
  assign _GEN_0_0 = io_fn[3];
  assign _GEN_8_0 = _T_24 | _T_25;
  assign _GEN_2_0 = _T_16 == _T_17;
  assign _GEN_5_1 = io_fn == 4'h6;
  assign _GEN_10_1 = _T_142 | _T_143;
  assign _GEN_7_2 = io_fn == 4'h1;
  assign _GEN_1_4 = io_fn[1];
  assign _GEN_4_2 = io_fn == 4'h4;
  assign _GEN_3_5 = _T_24 | _T_25;
  assign _GEN_6_5 = io_fn == 4'h7;
endmodule
module CSRFile( // @[:Sodor3Stage.fir@1547.2]
  input         metaReset,
  input         clock, // @[:Sodor3Stage.fir@1548.4]
  input         reset, // @[:Sodor3Stage.fir@1549.4]
  input  [2:0]  io_rw_cmd, // @[:Sodor3Stage.fir@1550.4]
  output [31:0] io_rw_rdata, // @[:Sodor3Stage.fir@1550.4]
  input  [31:0] io_rw_wdata, // @[:Sodor3Stage.fir@1550.4]
  output        io_eret, // @[:Sodor3Stage.fir@1550.4]
  input  [11:0] io_decode_csr, // @[:Sodor3Stage.fir@1550.4]
  output        io_status_debug, // @[:Sodor3Stage.fir@1550.4]
  output [1:0]  io_status_prv, // @[:Sodor3Stage.fir@1550.4]
  output        io_status_sd, // @[:Sodor3Stage.fir@1550.4]
  output [7:0]  io_status_zero1, // @[:Sodor3Stage.fir@1550.4]
  output        io_status_tsr, // @[:Sodor3Stage.fir@1550.4]
  output        io_status_tw, // @[:Sodor3Stage.fir@1550.4]
  output        io_status_tvm, // @[:Sodor3Stage.fir@1550.4]
  output        io_status_mxr, // @[:Sodor3Stage.fir@1550.4]
  output        io_status_sum, // @[:Sodor3Stage.fir@1550.4]
  output        io_status_mprv, // @[:Sodor3Stage.fir@1550.4]
  output [1:0]  io_status_xs, // @[:Sodor3Stage.fir@1550.4]
  output [1:0]  io_status_fs, // @[:Sodor3Stage.fir@1550.4]
  output [1:0]  io_status_mpp, // @[:Sodor3Stage.fir@1550.4]
  output [1:0]  io_status_hpp, // @[:Sodor3Stage.fir@1550.4]
  output        io_status_spp, // @[:Sodor3Stage.fir@1550.4]
  output        io_status_mpie, // @[:Sodor3Stage.fir@1550.4]
  output        io_status_hpie, // @[:Sodor3Stage.fir@1550.4]
  output        io_status_spie, // @[:Sodor3Stage.fir@1550.4]
  output        io_status_upie, // @[:Sodor3Stage.fir@1550.4]
  output        io_status_mie, // @[:Sodor3Stage.fir@1550.4]
  output        io_status_hie, // @[:Sodor3Stage.fir@1550.4]
  output        io_status_sie, // @[:Sodor3Stage.fir@1550.4]
  output        io_status_uie, // @[:Sodor3Stage.fir@1550.4]
  output [31:0] io_evec, // @[:Sodor3Stage.fir@1550.4]
  input         io_exception, // @[:Sodor3Stage.fir@1550.4]
  input         io_retire, // @[:Sodor3Stage.fir@1550.4]
  input  [31:0] io_pc, // @[:Sodor3Stage.fir@1550.4]
  output        _GEN_338_0,
  output        _GEN_224_0,
  output        _GEN_218_0,
  output        _GEN_323_0,
  output        _GEN_302_0,
  output        _GEN_239_0,
  output        _GEN_317_0,
  output        _GEN_385_0,
  output        _GEN_197_0,
  output        _GEN_296_0,
  output        _GEN_203_0,
  output        _GEN_212_0,
  output        _GEN_320_0,
  output        _GEN_200_0,
  output        _GEN_388_0,
  output        _GEN_191_0,
  output        _GEN_181_0,
  output        _GEN_190_1,
  output        _GEN_289_0,
  output        _GEN_299_0,
  output        _GEN_311_0,
  output        _GEN_206_0,
  output        _GEN_367_0,
  output        _GEN_175_0,
  output        _GEN_305_0,
  output        _GEN_274_0,
  output        _GEN_373_0,
  output        _GEN_376_0,
  output        _GEN_382_0,
  output        _GEN_370_0,
  output        _GEN_349_0,
  output        _GEN_262_0,
  output        _GEN_355_0,
  output        _GEN_277_0,
  output        _GEN_194_0,
  output        _GEN_184_0,
  output        _GEN_293_0,
  output        _GEN_157_0,
  output        _GEN_361_0,
  output        _GEN_256_0,
  output        _GEN_283_0,
  output        _GEN_163_0,
  output        _GEN_178_0,
  output        _GEN_11_0,
  output        _GEN_259_0,
  output        _GEN_358_0,
  output        _GEN_172_0,
  output        _GEN_271_0,
  output        _GEN_265_0,
  output        _GEN_280_0,
  output        _GEN_160_0,
  output        _GEN_343_0,
  output        _GEN_379_0,
  output        _GEN_238_0,
  output        _GEN_337_0,
  output        _GEN_364_0,
  output        _GEN_244_0,
  output        _GEN_166_0,
  output        _GEN_286_0,
  output        _GEN_151_0,
  output        _GEN_187_0,
  output        _GEN_319_1,
  output        _GEN_268_0,
  output        _GEN_226_1,
  output        _GEN_147_1,
  output        _GEN_352_0,
  output        _GEN_247_1,
  output        _GEN_325_1,
  output        _GEN_169_0,
  output        _GEN_232_1,
  output        _GEN_331_1,
  output        _GEN_346_0,
  output        _GEN_154_0,
  output        _GEN_340_0,
  output        _GEN_253_0,
  output        _GEN_211_1,
  output        _GEN_220_1,
  output        _GEN_229_1,
  output        _GEN_292_1,
  output        _GEN_307_1,
  output        _GEN_193_1,
  output        _GEN_313_1,
  output        _GEN_328_0,
  output        _GEN_235_0,
  output        _GEN_3_3,
  output        _GEN_250_0,
  output        _GEN_208_1,
  output        _GEN_214_1,
  output        _GEN_241_0,
  output        _GEN_334_0,
  output        _GEN_217_0,
  output        _GEN_316_0,
  output        _GEN_180_1,
  output        _GEN_384_1,
  output        _GEN_301_1,
  output        _GEN_196_1,
  output        _GEN_186_1,
  output        _GEN_295_1,
  output        _GEN_223_0,
  output        _GEN_322_0,
  output        _GEN_279_1,
  output        _GEN_310_1,
  output        _GEN_285_1,
  output        _GEN_202_1,
  output        _GEN_378_1,
  output        _GEN_351_1,
  output        _GEN_387_1,
  output        _GEN_189_1,
  output        _GEN_372_1,
  output        _GEN_267_1,
  output        _GEN_174_1,
  output        _GEN_205_1,
  output        _GEN_273_1,
  output        _GEN_168_1,
  output        _GEN_199_1,
  output        _GEN_298_1,
  output        _GEN_304_1,
  output        _GEN_366_1,
  output        _GEN_360_1,
  output        _GEN_288_1,
  output        _GEN_375_1,
  output        _GEN_255_1,
  output        _GEN_261_1,
  output        _GEN_270_1,
  output        _GEN_150_1,
  output        _GEN_333_1,
  output        _GEN_177_1,
  output        _GEN_381_1,
  output        _GEN_276_1,
  output        _GEN_354_1,
  output        _GEN_348_1,
  output        _GEN_249_1,
  output        _GEN_369_1,
  output        _GEN_183_1,
  output        _GEN_282_1,
  output        _GEN_162_1,
  output        _GEN_156_1,
  output        _GEN_165_1,
  output        _GEN_342_1,
  output        _GEN_264_1,
  output        _GEN_159_1,
  output        _GEN_222_1,
  output        _GEN_363_1,
  output        _GEN_357_1,
  output        _GEN_321_1,
  output        _GEN_7_3,
  output        _GEN_330_1,
  output        _GEN_243_1,
  output        _GEN_237_1,
  output        _GEN_315_1,
  output        _GEN_336_1,
  output        _GEN_258_1,
  output        _GEN_171_1,
  output        _GEN_303_1,
  output        _GEN_146_1,
  output        _GEN_225_1,
  output        _GEN_231_1,
  output        _GEN_240_1,
  output        _GEN_339_1,
  output        _GEN_153_1,
  output        _GEN_252_1,
  output        _GEN_297_1,
  output        _GEN_324_1,
  output        _GEN_219_1,
  output        _GEN_246_1,
  output        _GEN_318_1,
  output        _GEN_345_1,
  output        _GEN_204_1,
  output        _GEN_213_1,
  output        _GEN_228_1,
  output        _GEN_281_1,
  output        _GEN_234_1,
  output        _GEN_312_1,
  output        _GEN_192_1,
  output        _GEN_306_1,
  output        _GEN_207_1,
  output        _GEN_300_1,
  output        _GEN_327_1,
  output        _GEN_182_1,
  output        _GEN_291_1,
  output        _GEN_290_0,
  output        _GEN_383_1,
  output        _GEN_195_1,
  output        _GEN_185_1,
  output        _GEN_179_1,
  output        _GEN_216_1,
  output        _GEN_278_1,
  output        _GEN_201_1,
  output        _GEN_210_1,
  output        _GEN_263_1,
  output        _GEN_309_1,
  output        _GEN_164_1,
  output        _GEN_362_1,
  output        _GEN_377_1,
  output        _GEN_294_1,
  output        _GEN_284_1,
  output        _GEN_371_1,
  output        _GEN_260_1,
  output        _GEN_266_1,
  output        _GEN_380_1,
  output        _GEN_365_1,
  output        _GEN_251_1,
  output        _GEN_15_2,
  output        _GEN_359_1,
  output        _GEN_152_1,
  output        _GEN_188_1,
  output        _GEN_173_1,
  output        _GEN_287_1,
  output        _GEN_386_1,
  output        _GEN_245_1,
  output        _GEN_272_1,
  output        _GEN_344_1,
  output        _GEN_198_1,
  output        _GEN_167_1,
  output        _GEN_254_1,
  output        _GEN_161_1,
  output        _GEN_347_1,
  output        _GEN_170_1,
  output        _GEN_275_1,
  output        _GEN_269_1,
  output        _GEN_155_1,
  output        _GEN_368_1,
  output        _GEN_233_1,
  output        _GEN_227_1,
  output        _GEN_326_1,
  output        _GEN_149_1,
  output        _GEN_353_1,
  output        _GEN_248_1,
  output        _GEN_374_1,
  output        _GEN_332_1,
  output        _GEN_176_1,
  output        _GEN_314_1,
  output        _GEN_308_1,
  output        _GEN_341_1,
  output        _GEN_5_5,
  output        _GEN_356_1,
  output        _GEN_158_1,
  output        _GEN_209_1,
  output        _GEN_221_1,
  output        _GEN_236_1,
  output        _GEN_335_1,
  output        _GEN_329_1,
  output        _GEN_230_1,
  output        _GEN_242_1,
  output        _GEN_257_1,
  output        _GEN_350_1,
  output        _GEN_215_1
);
  reg [1:0] reg_mstatus_prv; // @[csr.scala 163:24:Sodor3Stage.fir@1726.4]
  reg [31:0] _RAND_0;
  reg  reg_mstatus_mpie; // @[csr.scala 163:24:Sodor3Stage.fir@1726.4]
  reg [31:0] _RAND_1;
  reg  reg_mstatus_mie; // @[csr.scala 163:24:Sodor3Stage.fir@1726.4]
  reg [31:0] _RAND_2;
  reg [31:0] reg_mepc; // @[csr.scala 164:21:Sodor3Stage.fir@1727.4]
  reg [31:0] _RAND_3;
  reg [31:0] reg_mcause; // @[csr.scala 165:23:Sodor3Stage.fir@1728.4]
  reg [31:0] _RAND_4;
  reg [31:0] reg_mtval; // @[csr.scala 166:22:Sodor3Stage.fir@1729.4]
  reg [31:0] _RAND_5;
  reg [31:0] reg_mscratch; // @[csr.scala 167:25:Sodor3Stage.fir@1730.4]
  reg [31:0] _RAND_6;
  reg [31:0] reg_medeleg; // @[csr.scala 169:24:Sodor3Stage.fir@1732.4]
  reg [31:0] _RAND_7;
  reg  reg_mip_mtip; // @[csr.scala 171:20:Sodor3Stage.fir@1768.4]
  reg [31:0] _RAND_8;
  reg  reg_mip_msip; // @[csr.scala 171:20:Sodor3Stage.fir@1768.4]
  reg [31:0] _RAND_9;
  reg  reg_mie_mtip; // @[csr.scala 172:20:Sodor3Stage.fir@1804.4]
  reg [31:0] _RAND_10;
  reg  reg_mie_msip; // @[csr.scala 172:20:Sodor3Stage.fir@1804.4]
  reg [31:0] _RAND_11;
  reg [5:0] _T_176; // @[util.scala 114:37:Sodor3Stage.fir@1807.4]
  reg [31:0] _RAND_12;
  reg [57:0] _T_180; // @[util.scala 119:27:Sodor3Stage.fir@1810.4]
  reg [63:0] _RAND_13;
  reg [5:0] _T_188; // @[util.scala 114:37:Sodor3Stage.fir@1818.4]
  reg [31:0] _RAND_14;
  reg [57:0] _T_192; // @[util.scala 119:27:Sodor3Stage.fir@1821.4]
  reg [63:0] _RAND_15;
  reg [39:0] _T_200; // @[util.scala 114:75:Sodor3Stage.fir@1830.4]
  reg [63:0] _RAND_16;
  reg [39:0] _T_203; // @[util.scala 114:75:Sodor3Stage.fir@1833.4]
  reg [63:0] _RAND_17;
  reg [39:0] _T_206; // @[util.scala 114:75:Sodor3Stage.fir@1836.4]
  reg [63:0] _RAND_18;
  reg [39:0] _T_209; // @[util.scala 114:75:Sodor3Stage.fir@1839.4]
  reg [63:0] _RAND_19;
  reg [39:0] _T_212; // @[util.scala 114:75:Sodor3Stage.fir@1842.4]
  reg [63:0] _RAND_20;
  reg [39:0] _T_215; // @[util.scala 114:75:Sodor3Stage.fir@1845.4]
  reg [63:0] _RAND_21;
  reg [39:0] _T_218; // @[util.scala 114:75:Sodor3Stage.fir@1848.4]
  reg [63:0] _RAND_22;
  reg [39:0] _T_221; // @[util.scala 114:75:Sodor3Stage.fir@1851.4]
  reg [63:0] _RAND_23;
  reg [39:0] _T_224; // @[util.scala 114:75:Sodor3Stage.fir@1854.4]
  reg [63:0] _RAND_24;
  reg [39:0] _T_227; // @[util.scala 114:75:Sodor3Stage.fir@1857.4]
  reg [63:0] _RAND_25;
  reg [39:0] _T_230; // @[util.scala 114:75:Sodor3Stage.fir@1860.4]
  reg [63:0] _RAND_26;
  reg [39:0] _T_233; // @[util.scala 114:75:Sodor3Stage.fir@1863.4]
  reg [63:0] _RAND_27;
  reg [39:0] _T_236; // @[util.scala 114:75:Sodor3Stage.fir@1866.4]
  reg [63:0] _RAND_28;
  reg [39:0] _T_239; // @[util.scala 114:75:Sodor3Stage.fir@1869.4]
  reg [63:0] _RAND_29;
  reg [39:0] _T_242; // @[util.scala 114:75:Sodor3Stage.fir@1872.4]
  reg [63:0] _RAND_30;
  reg [39:0] _T_245; // @[util.scala 114:75:Sodor3Stage.fir@1875.4]
  reg [63:0] _RAND_31;
  reg [39:0] _T_248; // @[util.scala 114:75:Sodor3Stage.fir@1878.4]
  reg [63:0] _RAND_32;
  reg [39:0] _T_251; // @[util.scala 114:75:Sodor3Stage.fir@1881.4]
  reg [63:0] _RAND_33;
  reg [39:0] _T_254; // @[util.scala 114:75:Sodor3Stage.fir@1884.4]
  reg [63:0] _RAND_34;
  reg [39:0] _T_257; // @[util.scala 114:75:Sodor3Stage.fir@1887.4]
  reg [63:0] _RAND_35;
  reg [39:0] _T_260; // @[util.scala 114:75:Sodor3Stage.fir@1890.4]
  reg [63:0] _RAND_36;
  reg [39:0] _T_263; // @[util.scala 114:75:Sodor3Stage.fir@1893.4]
  reg [63:0] _RAND_37;
  reg [39:0] _T_266; // @[util.scala 114:75:Sodor3Stage.fir@1896.4]
  reg [63:0] _RAND_38;
  reg [39:0] _T_269; // @[util.scala 114:75:Sodor3Stage.fir@1899.4]
  reg [63:0] _RAND_39;
  reg [39:0] _T_272; // @[util.scala 114:75:Sodor3Stage.fir@1902.4]
  reg [63:0] _RAND_40;
  reg [39:0] _T_275; // @[util.scala 114:75:Sodor3Stage.fir@1905.4]
  reg [63:0] _RAND_41;
  reg [39:0] _T_278; // @[util.scala 114:75:Sodor3Stage.fir@1908.4]
  reg [63:0] _RAND_42;
  reg [39:0] _T_281; // @[util.scala 114:75:Sodor3Stage.fir@1911.4]
  reg [63:0] _RAND_43;
  reg [39:0] _T_284; // @[util.scala 114:75:Sodor3Stage.fir@1914.4]
  reg [63:0] _RAND_44;
  reg [39:0] _T_287; // @[util.scala 114:75:Sodor3Stage.fir@1917.4]
  reg [63:0] _RAND_45;
  reg [39:0] _T_290; // @[util.scala 114:75:Sodor3Stage.fir@1920.4]
  reg [63:0] _RAND_46;
  reg [39:0] _T_293; // @[util.scala 114:75:Sodor3Stage.fir@1923.4]
  reg [63:0] _RAND_47;
  reg [31:0] reg_dpc; // @[csr.scala 188:20:Sodor3Stage.fir@2014.4]
  reg [31:0] _RAND_48;
  reg [31:0] reg_dscratch; // @[csr.scala 189:25:Sodor3Stage.fir@2015.4]
  reg [31:0] _RAND_49;
  reg  reg_dcsr_ebreakm; // @[csr.scala 194:21:Sodor3Stage.fir@2068.4]
  reg [31:0] _RAND_50;
  reg  reg_dcsr_step; // @[csr.scala 194:21:Sodor3Stage.fir@2068.4]
  reg [31:0] _RAND_51;
  wire [6:0] _T_177; // @[util.scala 115:33:Sodor3Stage.fir@1808.4]
  wire  _T_181; // @[util.scala 120:20:Sodor3Stage.fir@1811.4]
  wire [58:0] _T_183; // @[util.scala 120:43:Sodor3Stage.fir@1813.6]
  wire [57:0] _T_184; // @[util.scala 120:43:Sodor3Stage.fir@1814.6]
  wire [63:0] _T_185; // @[Cat.scala 30:58:Sodor3Stage.fir@1817.4]
  wire [5:0] _GEN_389; // @[util.scala 115:33:Sodor3Stage.fir@1819.4]
  wire [6:0] _T_189; // @[util.scala 115:33:Sodor3Stage.fir@1819.4]
  wire  _T_193; // @[util.scala 120:20:Sodor3Stage.fir@1822.4]
  wire [58:0] _T_195; // @[util.scala 120:43:Sodor3Stage.fir@1824.6]
  wire [57:0] _T_196; // @[util.scala 120:43:Sodor3Stage.fir@1825.6]
  wire [63:0] _T_197; // @[Cat.scala 30:58:Sodor3Stage.fir@1828.4]
  wire [40:0] _T_201; // @[util.scala 115:33:Sodor3Stage.fir@1831.4]
  wire [40:0] _T_204; // @[util.scala 115:33:Sodor3Stage.fir@1834.4]
  wire [40:0] _T_207; // @[util.scala 115:33:Sodor3Stage.fir@1837.4]
  wire [40:0] _T_210; // @[util.scala 115:33:Sodor3Stage.fir@1840.4]
  wire [40:0] _T_213; // @[util.scala 115:33:Sodor3Stage.fir@1843.4]
  wire [40:0] _T_216; // @[util.scala 115:33:Sodor3Stage.fir@1846.4]
  wire [40:0] _T_219; // @[util.scala 115:33:Sodor3Stage.fir@1849.4]
  wire [40:0] _T_222; // @[util.scala 115:33:Sodor3Stage.fir@1852.4]
  wire [40:0] _T_225; // @[util.scala 115:33:Sodor3Stage.fir@1855.4]
  wire [40:0] _T_228; // @[util.scala 115:33:Sodor3Stage.fir@1858.4]
  wire [40:0] _T_231; // @[util.scala 115:33:Sodor3Stage.fir@1861.4]
  wire [40:0] _T_234; // @[util.scala 115:33:Sodor3Stage.fir@1864.4]
  wire [40:0] _T_237; // @[util.scala 115:33:Sodor3Stage.fir@1867.4]
  wire [40:0] _T_240; // @[util.scala 115:33:Sodor3Stage.fir@1870.4]
  wire [40:0] _T_243; // @[util.scala 115:33:Sodor3Stage.fir@1873.4]
  wire [40:0] _T_246; // @[util.scala 115:33:Sodor3Stage.fir@1876.4]
  wire [40:0] _T_249; // @[util.scala 115:33:Sodor3Stage.fir@1879.4]
  wire [40:0] _T_252; // @[util.scala 115:33:Sodor3Stage.fir@1882.4]
  wire [40:0] _T_255; // @[util.scala 115:33:Sodor3Stage.fir@1885.4]
  wire [40:0] _T_258; // @[util.scala 115:33:Sodor3Stage.fir@1888.4]
  wire [40:0] _T_261; // @[util.scala 115:33:Sodor3Stage.fir@1891.4]
  wire [40:0] _T_264; // @[util.scala 115:33:Sodor3Stage.fir@1894.4]
  wire [40:0] _T_267; // @[util.scala 115:33:Sodor3Stage.fir@1897.4]
  wire [40:0] _T_270; // @[util.scala 115:33:Sodor3Stage.fir@1900.4]
  wire [40:0] _T_273; // @[util.scala 115:33:Sodor3Stage.fir@1903.4]
  wire [40:0] _T_276; // @[util.scala 115:33:Sodor3Stage.fir@1906.4]
  wire [40:0] _T_279; // @[util.scala 115:33:Sodor3Stage.fir@1909.4]
  wire [40:0] _T_282; // @[util.scala 115:33:Sodor3Stage.fir@1912.4]
  wire [40:0] _T_285; // @[util.scala 115:33:Sodor3Stage.fir@1915.4]
  wire [40:0] _T_288; // @[util.scala 115:33:Sodor3Stage.fir@1918.4]
  wire [40:0] _T_291; // @[util.scala 115:33:Sodor3Stage.fir@1921.4]
  wire [40:0] _T_294; // @[util.scala 115:33:Sodor3Stage.fir@1924.4]
  wire  system_insn; // @[csr.scala 196:31:Sodor3Stage.fir@2069.4]
  wire  _T_410; // @[csr.scala 197:27:Sodor3Stage.fir@2070.4]
  wire  _T_412; // @[csr.scala 197:39:Sodor3Stage.fir@2071.4]
  wire  cpu_ren; // @[csr.scala 197:36:Sodor3Stage.fir@2072.4]
  wire [1:0] _T_413; // @[:Sodor3Stage.fir@2073.4]
  wire [1:0] _T_414; // @[:Sodor3Stage.fir@2074.4]
  wire [2:0] _T_415; // @[:Sodor3Stage.fir@2075.4]
  wire [4:0] _T_416; // @[:Sodor3Stage.fir@2076.4]
  wire [1:0] _T_417; // @[:Sodor3Stage.fir@2077.4]
  wire [2:0] _T_418; // @[:Sodor3Stage.fir@2078.4]
  wire [3:0] _T_419; // @[:Sodor3Stage.fir@2079.4]
  wire [4:0] _T_420; // @[:Sodor3Stage.fir@2080.4]
  wire [7:0] _T_421; // @[:Sodor3Stage.fir@2081.4]
  wire [12:0] _T_422; // @[:Sodor3Stage.fir@2082.4]
  wire [2:0] _T_423; // @[:Sodor3Stage.fir@2083.4]
  wire [4:0] _T_424; // @[:Sodor3Stage.fir@2084.4]
  wire [1:0] _T_425; // @[:Sodor3Stage.fir@2085.4]
  wire [2:0] _T_426; // @[:Sodor3Stage.fir@2086.4]
  wire [7:0] _T_427; // @[:Sodor3Stage.fir@2087.4]
  wire [8:0] _T_428; // @[:Sodor3Stage.fir@2088.4]
  wire [9:0] _T_429; // @[:Sodor3Stage.fir@2089.4]
  wire [2:0] _T_430; // @[:Sodor3Stage.fir@2090.4]
  wire [3:0] _T_431; // @[:Sodor3Stage.fir@2091.4]
  wire [13:0] _T_432; // @[:Sodor3Stage.fir@2092.4]
  wire [21:0] _T_433; // @[:Sodor3Stage.fir@2093.4]
  wire [34:0] read_mstatus; // @[:Sodor3Stage.fir@2094.4]
  wire [1:0] _T_441; // @[:Sodor3Stage.fir@2096.4]
  wire [3:0] _T_442; // @[:Sodor3Stage.fir@2097.4]
  wire [1:0] _T_444; // @[:Sodor3Stage.fir@2099.4]
  wire [3:0] _T_445; // @[:Sodor3Stage.fir@2100.4]
  wire [7:0] _T_446; // @[:Sodor3Stage.fir@2101.4]
  wire [15:0] _T_454; // @[:Sodor3Stage.fir@2109.4]
  wire [1:0] _T_456; // @[:Sodor3Stage.fir@2111.4]
  wire [3:0] _T_457; // @[:Sodor3Stage.fir@2112.4]
  wire [1:0] _T_459; // @[:Sodor3Stage.fir@2114.4]
  wire [3:0] _T_460; // @[:Sodor3Stage.fir@2115.4]
  wire [7:0] _T_461; // @[:Sodor3Stage.fir@2116.4]
  wire [15:0] _T_469; // @[:Sodor3Stage.fir@2124.4]
  wire [2:0] _T_470; // @[csr.scala 222:27:Sodor3Stage.fir@2125.4]
  wire [4:0] _T_471; // @[csr.scala 222:27:Sodor3Stage.fir@2126.4]
  wire [10:0] _T_475; // @[csr.scala 222:27:Sodor3Stage.fir@2130.4]
  wire [12:0] _T_479; // @[csr.scala 222:27:Sodor3Stage.fir@2134.4]
  wire [16:0] _T_481; // @[csr.scala 222:27:Sodor3Stage.fir@2136.4]
  wire [20:0] _T_482; // @[csr.scala 222:27:Sodor3Stage.fir@2137.4]
  wire [31:0] _T_483; // @[csr.scala 222:27:Sodor3Stage.fir@2138.4]
  wire  _T_487; // @[csr.scala 259:76:Sodor3Stage.fir@2139.4]
  wire  _T_489; // @[csr.scala 259:76:Sodor3Stage.fir@2140.4]
  wire  _T_491; // @[csr.scala 259:76:Sodor3Stage.fir@2141.4]
  wire  _T_497; // @[csr.scala 259:76:Sodor3Stage.fir@2144.4]
  wire  _T_499; // @[csr.scala 259:76:Sodor3Stage.fir@2145.4]
  wire  _T_501; // @[csr.scala 259:76:Sodor3Stage.fir@2146.4]
  wire  _T_503; // @[csr.scala 259:76:Sodor3Stage.fir@2147.4]
  wire  _T_505; // @[csr.scala 259:76:Sodor3Stage.fir@2148.4]
  wire  _T_507; // @[csr.scala 259:76:Sodor3Stage.fir@2149.4]
  wire  _T_509; // @[csr.scala 259:76:Sodor3Stage.fir@2150.4]
  wire  _T_511; // @[csr.scala 259:76:Sodor3Stage.fir@2151.4]
  wire  _T_513; // @[csr.scala 259:76:Sodor3Stage.fir@2152.4]
  wire  _T_517; // @[csr.scala 259:76:Sodor3Stage.fir@2154.4]
  wire  _T_519; // @[csr.scala 259:76:Sodor3Stage.fir@2155.4]
  wire  _T_521; // @[csr.scala 259:76:Sodor3Stage.fir@2156.4]
  wire  _T_523; // @[csr.scala 259:76:Sodor3Stage.fir@2157.4]
  wire  _T_525; // @[csr.scala 259:76:Sodor3Stage.fir@2158.4]
  wire  _T_527; // @[csr.scala 259:76:Sodor3Stage.fir@2159.4]
  wire  _T_529; // @[csr.scala 259:76:Sodor3Stage.fir@2160.4]
  wire  _T_531; // @[csr.scala 259:76:Sodor3Stage.fir@2161.4]
  wire  _T_533; // @[csr.scala 259:76:Sodor3Stage.fir@2162.4]
  wire  _T_535; // @[csr.scala 259:76:Sodor3Stage.fir@2163.4]
  wire  _T_537; // @[csr.scala 259:76:Sodor3Stage.fir@2164.4]
  wire  _T_539; // @[csr.scala 259:76:Sodor3Stage.fir@2165.4]
  wire  _T_541; // @[csr.scala 259:76:Sodor3Stage.fir@2166.4]
  wire  _T_543; // @[csr.scala 259:76:Sodor3Stage.fir@2167.4]
  wire  _T_545; // @[csr.scala 259:76:Sodor3Stage.fir@2168.4]
  wire  _T_547; // @[csr.scala 259:76:Sodor3Stage.fir@2169.4]
  wire  _T_549; // @[csr.scala 259:76:Sodor3Stage.fir@2170.4]
  wire  _T_551; // @[csr.scala 259:76:Sodor3Stage.fir@2171.4]
  wire  _T_553; // @[csr.scala 259:76:Sodor3Stage.fir@2172.4]
  wire  _T_555; // @[csr.scala 259:76:Sodor3Stage.fir@2173.4]
  wire  _T_557; // @[csr.scala 259:76:Sodor3Stage.fir@2174.4]
  wire  _T_559; // @[csr.scala 259:76:Sodor3Stage.fir@2175.4]
  wire  _T_561; // @[csr.scala 259:76:Sodor3Stage.fir@2176.4]
  wire  _T_563; // @[csr.scala 259:76:Sodor3Stage.fir@2177.4]
  wire  _T_565; // @[csr.scala 259:76:Sodor3Stage.fir@2178.4]
  wire  _T_567; // @[csr.scala 259:76:Sodor3Stage.fir@2179.4]
  wire  _T_569; // @[csr.scala 259:76:Sodor3Stage.fir@2180.4]
  wire  _T_571; // @[csr.scala 259:76:Sodor3Stage.fir@2181.4]
  wire  _T_573; // @[csr.scala 259:76:Sodor3Stage.fir@2182.4]
  wire  _T_575; // @[csr.scala 259:76:Sodor3Stage.fir@2183.4]
  wire  _T_577; // @[csr.scala 259:76:Sodor3Stage.fir@2184.4]
  wire  _T_579; // @[csr.scala 259:76:Sodor3Stage.fir@2185.4]
  wire  _T_581; // @[csr.scala 259:76:Sodor3Stage.fir@2186.4]
  wire  _T_583; // @[csr.scala 259:76:Sodor3Stage.fir@2187.4]
  wire  _T_585; // @[csr.scala 259:76:Sodor3Stage.fir@2188.4]
  wire  _T_587; // @[csr.scala 259:76:Sodor3Stage.fir@2189.4]
  wire  _T_589; // @[csr.scala 259:76:Sodor3Stage.fir@2190.4]
  wire  _T_591; // @[csr.scala 259:76:Sodor3Stage.fir@2191.4]
  wire  _T_593; // @[csr.scala 259:76:Sodor3Stage.fir@2192.4]
  wire  _T_595; // @[csr.scala 259:76:Sodor3Stage.fir@2193.4]
  wire  _T_597; // @[csr.scala 259:76:Sodor3Stage.fir@2194.4]
  wire  _T_599; // @[csr.scala 259:76:Sodor3Stage.fir@2195.4]
  wire  _T_601; // @[csr.scala 259:76:Sodor3Stage.fir@2196.4]
  wire  _T_603; // @[csr.scala 259:76:Sodor3Stage.fir@2197.4]
  wire  _T_605; // @[csr.scala 259:76:Sodor3Stage.fir@2198.4]
  wire  _T_607; // @[csr.scala 259:76:Sodor3Stage.fir@2199.4]
  wire  _T_609; // @[csr.scala 259:76:Sodor3Stage.fir@2200.4]
  wire  _T_611; // @[csr.scala 259:76:Sodor3Stage.fir@2201.4]
  wire  _T_613; // @[csr.scala 259:76:Sodor3Stage.fir@2202.4]
  wire  _T_615; // @[csr.scala 259:76:Sodor3Stage.fir@2203.4]
  wire  _T_617; // @[csr.scala 259:76:Sodor3Stage.fir@2204.4]
  wire  _T_619; // @[csr.scala 259:76:Sodor3Stage.fir@2205.4]
  wire  _T_621; // @[csr.scala 259:76:Sodor3Stage.fir@2206.4]
  wire  _T_623; // @[csr.scala 259:76:Sodor3Stage.fir@2207.4]
  wire  _T_625; // @[csr.scala 259:76:Sodor3Stage.fir@2208.4]
  wire  _T_627; // @[csr.scala 259:76:Sodor3Stage.fir@2209.4]
  wire  _T_629; // @[csr.scala 259:76:Sodor3Stage.fir@2210.4]
  wire  _T_631; // @[csr.scala 259:76:Sodor3Stage.fir@2211.4]
  wire  _T_633; // @[csr.scala 259:76:Sodor3Stage.fir@2212.4]
  wire  _T_635; // @[csr.scala 259:76:Sodor3Stage.fir@2213.4]
  wire  _T_637; // @[csr.scala 259:76:Sodor3Stage.fir@2214.4]
  wire  _T_639; // @[csr.scala 259:76:Sodor3Stage.fir@2215.4]
  wire  _T_641; // @[csr.scala 259:76:Sodor3Stage.fir@2216.4]
  wire  _T_643; // @[csr.scala 259:76:Sodor3Stage.fir@2217.4]
  wire  _T_645; // @[csr.scala 259:76:Sodor3Stage.fir@2218.4]
  wire  _T_647; // @[csr.scala 259:76:Sodor3Stage.fir@2219.4]
  wire  _T_649; // @[csr.scala 259:76:Sodor3Stage.fir@2220.4]
  wire  _T_651; // @[csr.scala 259:76:Sodor3Stage.fir@2221.4]
  wire  _T_653; // @[csr.scala 259:76:Sodor3Stage.fir@2222.4]
  wire  _T_655; // @[csr.scala 259:76:Sodor3Stage.fir@2223.4]
  wire [1:0] _T_656; // @[csr.scala 261:57:Sodor3Stage.fir@2224.4]
  wire  priv_sufficient; // @[csr.scala 261:41:Sodor3Stage.fir@2225.4]
  wire [1:0] _T_657; // @[csr.scala 262:32:Sodor3Stage.fir@2226.4]
  wire [1:0] _T_658; // @[csr.scala 262:40:Sodor3Stage.fir@2227.4]
  wire  read_only; // @[csr.scala 262:40:Sodor3Stage.fir@2228.4]
  wire  _T_660; // @[csr.scala 263:38:Sodor3Stage.fir@2229.4]
  wire  _T_661; // @[csr.scala 263:25:Sodor3Stage.fir@2230.4]
  wire  cpu_wen; // @[csr.scala 263:47:Sodor3Stage.fir@2231.4]
  wire  _T_663; // @[csr.scala 264:24:Sodor3Stage.fir@2232.4]
  wire  wen; // @[csr.scala 264:21:Sodor3Stage.fir@2233.4]
  wire  _T_664; // @[util.scala 25:47:Sodor3Stage.fir@2234.4]
  wire  _T_665; // @[util.scala 25:47:Sodor3Stage.fir@2235.4]
  wire  _T_666; // @[util.scala 25:62:Sodor3Stage.fir@2236.4]
  wire [31:0] _T_668; // @[csr.scala 390:9:Sodor3Stage.fir@2237.4]
  wire [31:0] _T_669; // @[csr.scala 390:53:Sodor3Stage.fir@2238.4]
  wire [31:0] _T_672; // @[csr.scala 390:68:Sodor3Stage.fir@2240.4]
  wire [31:0] _T_673; // @[csr.scala 390:64:Sodor3Stage.fir@2241.4]
  wire [31:0] wdata; // @[csr.scala 390:62:Sodor3Stage.fir@2242.4]
  wire [2:0] _T_675; // @[csr.scala 267:36:Sodor3Stage.fir@2243.4]
  wire [7:0] opcode; // @[csr.scala 267:20:Sodor3Stage.fir@2244.4]
  wire  _T_676; // @[csr.scala 268:40:Sodor3Stage.fir@2245.4]
  wire  insn_call; // @[csr.scala 268:31:Sodor3Stage.fir@2246.4]
  wire  _T_677; // @[csr.scala 269:41:Sodor3Stage.fir@2247.4]
  wire  insn_break; // @[csr.scala 269:32:Sodor3Stage.fir@2248.4]
  wire  _T_678; // @[csr.scala 270:39:Sodor3Stage.fir@2249.4]
  wire  _T_679; // @[csr.scala 270:30:Sodor3Stage.fir@2250.4]
  wire  insn_ret; // @[csr.scala 270:43:Sodor3Stage.fir@2251.4]
  wire  _T_962; // @[csr.scala 282:24:Sodor3Stage.fir@2469.4]
  wire [31:0] _GEN_4; // @[csr.scala 285:23:Sodor3Stage.fir@2472.4]
  wire [1:0] _T_966; // @[Bitwise.scala 48:55:Sodor3Stage.fir@2477.4]
  wire  _T_968; // @[csr.scala 291:52:Sodor3Stage.fir@2478.4]
  wire  _T_970; // @[csr.scala 291:9:Sodor3Stage.fir@2480.4]
  wire  _T_975; // @[csr.scala 298:33:Sodor3Stage.fir@2490.4]
  wire  _T_976; // @[csr.scala 298:17:Sodor3Stage.fir@2491.4]
  wire [31:0] _GEN_8; // @[csr.scala 298:38:Sodor3Stage.fir@2492.4]
  wire  _T_980; // @[csr.scala 305:21:Sodor3Stage.fir@2498.4]
  wire  _T_981; // @[csr.scala 305:18:Sodor3Stage.fir@2499.4]
  wire [31:0] _GEN_12; // @[csr.scala 305:41:Sodor3Stage.fir@2500.4]
  wire [3:0] _GEN_390; // @[csr.scala 315:35:Sodor3Stage.fir@2508.6]
  wire [4:0] _T_985; // @[csr.scala 315:35:Sodor3Stage.fir@2508.6]
  wire [3:0] _T_986; // @[csr.scala 315:35:Sodor3Stage.fir@2509.6]
  wire [31:0] _GEN_13; // @[csr.scala 313:18:Sodor3Stage.fir@2506.4]
  wire [63:0] _T_991; // @[Mux.scala 19:72:Sodor3Stage.fir@2518.4]
  wire [63:0] _T_993; // @[Mux.scala 19:72:Sodor3Stage.fir@2519.4]
  wire [15:0] _T_995; // @[Mux.scala 19:72:Sodor3Stage.fir@2520.4]
  wire [8:0] _T_1001; // @[Mux.scala 19:72:Sodor3Stage.fir@2523.4]
  wire [34:0] _T_1003; // @[Mux.scala 19:72:Sodor3Stage.fir@2524.4]
  wire [8:0] _T_1005; // @[Mux.scala 19:72:Sodor3Stage.fir@2525.4]
  wire [15:0] _T_1007; // @[Mux.scala 19:72:Sodor3Stage.fir@2526.4]
  wire [15:0] _T_1009; // @[Mux.scala 19:72:Sodor3Stage.fir@2527.4]
  wire [31:0] _T_1011; // @[Mux.scala 19:72:Sodor3Stage.fir@2528.4]
  wire [31:0] _T_1013; // @[Mux.scala 19:72:Sodor3Stage.fir@2529.4]
  wire [31:0] _T_1015; // @[Mux.scala 19:72:Sodor3Stage.fir@2530.4]
  wire [31:0] _T_1017; // @[Mux.scala 19:72:Sodor3Stage.fir@2531.4]
  wire [31:0] _T_1021; // @[Mux.scala 19:72:Sodor3Stage.fir@2533.4]
  wire [31:0] _T_1023; // @[Mux.scala 19:72:Sodor3Stage.fir@2534.4]
  wire [31:0] _T_1025; // @[Mux.scala 19:72:Sodor3Stage.fir@2535.4]
  wire [31:0] _T_1027; // @[Mux.scala 19:72:Sodor3Stage.fir@2536.4]
  wire [39:0] _T_1029; // @[Mux.scala 19:72:Sodor3Stage.fir@2537.4]
  wire [39:0] _T_1031; // @[Mux.scala 19:72:Sodor3Stage.fir@2538.4]
  wire [39:0] _T_1033; // @[Mux.scala 19:72:Sodor3Stage.fir@2539.4]
  wire [39:0] _T_1035; // @[Mux.scala 19:72:Sodor3Stage.fir@2540.4]
  wire [39:0] _T_1037; // @[Mux.scala 19:72:Sodor3Stage.fir@2541.4]
  wire [39:0] _T_1039; // @[Mux.scala 19:72:Sodor3Stage.fir@2542.4]
  wire [39:0] _T_1041; // @[Mux.scala 19:72:Sodor3Stage.fir@2543.4]
  wire [39:0] _T_1043; // @[Mux.scala 19:72:Sodor3Stage.fir@2544.4]
  wire [39:0] _T_1045; // @[Mux.scala 19:72:Sodor3Stage.fir@2545.4]
  wire [39:0] _T_1047; // @[Mux.scala 19:72:Sodor3Stage.fir@2546.4]
  wire [39:0] _T_1049; // @[Mux.scala 19:72:Sodor3Stage.fir@2547.4]
  wire [39:0] _T_1051; // @[Mux.scala 19:72:Sodor3Stage.fir@2548.4]
  wire [39:0] _T_1053; // @[Mux.scala 19:72:Sodor3Stage.fir@2549.4]
  wire [39:0] _T_1055; // @[Mux.scala 19:72:Sodor3Stage.fir@2550.4]
  wire [39:0] _T_1057; // @[Mux.scala 19:72:Sodor3Stage.fir@2551.4]
  wire [39:0] _T_1059; // @[Mux.scala 19:72:Sodor3Stage.fir@2552.4]
  wire [39:0] _T_1061; // @[Mux.scala 19:72:Sodor3Stage.fir@2553.4]
  wire [39:0] _T_1063; // @[Mux.scala 19:72:Sodor3Stage.fir@2554.4]
  wire [39:0] _T_1065; // @[Mux.scala 19:72:Sodor3Stage.fir@2555.4]
  wire [39:0] _T_1067; // @[Mux.scala 19:72:Sodor3Stage.fir@2556.4]
  wire [39:0] _T_1069; // @[Mux.scala 19:72:Sodor3Stage.fir@2557.4]
  wire [39:0] _T_1071; // @[Mux.scala 19:72:Sodor3Stage.fir@2558.4]
  wire [39:0] _T_1073; // @[Mux.scala 19:72:Sodor3Stage.fir@2559.4]
  wire [39:0] _T_1075; // @[Mux.scala 19:72:Sodor3Stage.fir@2560.4]
  wire [39:0] _T_1077; // @[Mux.scala 19:72:Sodor3Stage.fir@2561.4]
  wire [39:0] _T_1079; // @[Mux.scala 19:72:Sodor3Stage.fir@2562.4]
  wire [39:0] _T_1081; // @[Mux.scala 19:72:Sodor3Stage.fir@2563.4]
  wire [39:0] _T_1083; // @[Mux.scala 19:72:Sodor3Stage.fir@2564.4]
  wire [39:0] _T_1085; // @[Mux.scala 19:72:Sodor3Stage.fir@2565.4]
  wire [39:0] _T_1087; // @[Mux.scala 19:72:Sodor3Stage.fir@2566.4]
  wire [39:0] _T_1089; // @[Mux.scala 19:72:Sodor3Stage.fir@2567.4]
  wire [39:0] _T_1091; // @[Mux.scala 19:72:Sodor3Stage.fir@2568.4]
  wire [39:0] _T_1093; // @[Mux.scala 19:72:Sodor3Stage.fir@2569.4]
  wire [39:0] _T_1095; // @[Mux.scala 19:72:Sodor3Stage.fir@2570.4]
  wire [39:0] _T_1097; // @[Mux.scala 19:72:Sodor3Stage.fir@2571.4]
  wire [39:0] _T_1099; // @[Mux.scala 19:72:Sodor3Stage.fir@2572.4]
  wire [39:0] _T_1101; // @[Mux.scala 19:72:Sodor3Stage.fir@2573.4]
  wire [39:0] _T_1103; // @[Mux.scala 19:72:Sodor3Stage.fir@2574.4]
  wire [39:0] _T_1105; // @[Mux.scala 19:72:Sodor3Stage.fir@2575.4]
  wire [39:0] _T_1107; // @[Mux.scala 19:72:Sodor3Stage.fir@2576.4]
  wire [39:0] _T_1109; // @[Mux.scala 19:72:Sodor3Stage.fir@2577.4]
  wire [39:0] _T_1111; // @[Mux.scala 19:72:Sodor3Stage.fir@2578.4]
  wire [39:0] _T_1113; // @[Mux.scala 19:72:Sodor3Stage.fir@2579.4]
  wire [39:0] _T_1115; // @[Mux.scala 19:72:Sodor3Stage.fir@2580.4]
  wire [39:0] _T_1117; // @[Mux.scala 19:72:Sodor3Stage.fir@2581.4]
  wire [39:0] _T_1119; // @[Mux.scala 19:72:Sodor3Stage.fir@2582.4]
  wire [39:0] _T_1121; // @[Mux.scala 19:72:Sodor3Stage.fir@2583.4]
  wire [39:0] _T_1123; // @[Mux.scala 19:72:Sodor3Stage.fir@2584.4]
  wire [39:0] _T_1125; // @[Mux.scala 19:72:Sodor3Stage.fir@2585.4]
  wire [39:0] _T_1127; // @[Mux.scala 19:72:Sodor3Stage.fir@2586.4]
  wire [39:0] _T_1129; // @[Mux.scala 19:72:Sodor3Stage.fir@2587.4]
  wire [39:0] _T_1131; // @[Mux.scala 19:72:Sodor3Stage.fir@2588.4]
  wire [39:0] _T_1133; // @[Mux.scala 19:72:Sodor3Stage.fir@2589.4]
  wire [39:0] _T_1135; // @[Mux.scala 19:72:Sodor3Stage.fir@2590.4]
  wire [39:0] _T_1137; // @[Mux.scala 19:72:Sodor3Stage.fir@2591.4]
  wire [39:0] _T_1139; // @[Mux.scala 19:72:Sodor3Stage.fir@2592.4]
  wire [39:0] _T_1141; // @[Mux.scala 19:72:Sodor3Stage.fir@2593.4]
  wire [39:0] _T_1143; // @[Mux.scala 19:72:Sodor3Stage.fir@2594.4]
  wire [39:0] _T_1145; // @[Mux.scala 19:72:Sodor3Stage.fir@2595.4]
  wire [39:0] _T_1147; // @[Mux.scala 19:72:Sodor3Stage.fir@2596.4]
  wire [39:0] _T_1149; // @[Mux.scala 19:72:Sodor3Stage.fir@2597.4]
  wire [39:0] _T_1151; // @[Mux.scala 19:72:Sodor3Stage.fir@2598.4]
  wire [39:0] _T_1153; // @[Mux.scala 19:72:Sodor3Stage.fir@2599.4]
  wire [39:0] _T_1155; // @[Mux.scala 19:72:Sodor3Stage.fir@2600.4]
  wire [63:0] _T_1160; // @[Mux.scala 19:72:Sodor3Stage.fir@2603.4]
  wire [63:0] _GEN_391; // @[Mux.scala 19:72:Sodor3Stage.fir@2604.4]
  wire [63:0] _T_1161; // @[Mux.scala 19:72:Sodor3Stage.fir@2604.4]
  wire [63:0] _GEN_392; // @[Mux.scala 19:72:Sodor3Stage.fir@2607.4]
  wire [63:0] _T_1164; // @[Mux.scala 19:72:Sodor3Stage.fir@2607.4]
  wire [63:0] _GEN_393; // @[Mux.scala 19:72:Sodor3Stage.fir@2608.4]
  wire [63:0] _T_1165; // @[Mux.scala 19:72:Sodor3Stage.fir@2608.4]
  wire [63:0] _GEN_394; // @[Mux.scala 19:72:Sodor3Stage.fir@2609.4]
  wire [63:0] _T_1166; // @[Mux.scala 19:72:Sodor3Stage.fir@2609.4]
  wire [63:0] _GEN_395; // @[Mux.scala 19:72:Sodor3Stage.fir@2610.4]
  wire [63:0] _T_1167; // @[Mux.scala 19:72:Sodor3Stage.fir@2610.4]
  wire [63:0] _GEN_396; // @[Mux.scala 19:72:Sodor3Stage.fir@2611.4]
  wire [63:0] _T_1168; // @[Mux.scala 19:72:Sodor3Stage.fir@2611.4]
  wire [63:0] _GEN_397; // @[Mux.scala 19:72:Sodor3Stage.fir@2612.4]
  wire [63:0] _T_1169; // @[Mux.scala 19:72:Sodor3Stage.fir@2612.4]
  wire [63:0] _GEN_398; // @[Mux.scala 19:72:Sodor3Stage.fir@2613.4]
  wire [63:0] _T_1170; // @[Mux.scala 19:72:Sodor3Stage.fir@2613.4]
  wire [63:0] _GEN_399; // @[Mux.scala 19:72:Sodor3Stage.fir@2614.4]
  wire [63:0] _T_1171; // @[Mux.scala 19:72:Sodor3Stage.fir@2614.4]
  wire [63:0] _GEN_400; // @[Mux.scala 19:72:Sodor3Stage.fir@2615.4]
  wire [63:0] _T_1172; // @[Mux.scala 19:72:Sodor3Stage.fir@2615.4]
  wire [63:0] _GEN_401; // @[Mux.scala 19:72:Sodor3Stage.fir@2617.4]
  wire [63:0] _T_1174; // @[Mux.scala 19:72:Sodor3Stage.fir@2617.4]
  wire [63:0] _GEN_402; // @[Mux.scala 19:72:Sodor3Stage.fir@2618.4]
  wire [63:0] _T_1175; // @[Mux.scala 19:72:Sodor3Stage.fir@2618.4]
  wire [63:0] _GEN_403; // @[Mux.scala 19:72:Sodor3Stage.fir@2619.4]
  wire [63:0] _T_1176; // @[Mux.scala 19:72:Sodor3Stage.fir@2619.4]
  wire [63:0] _GEN_404; // @[Mux.scala 19:72:Sodor3Stage.fir@2620.4]
  wire [63:0] _T_1177; // @[Mux.scala 19:72:Sodor3Stage.fir@2620.4]
  wire [63:0] _GEN_405; // @[Mux.scala 19:72:Sodor3Stage.fir@2621.4]
  wire [63:0] _T_1178; // @[Mux.scala 19:72:Sodor3Stage.fir@2621.4]
  wire [63:0] _GEN_406; // @[Mux.scala 19:72:Sodor3Stage.fir@2622.4]
  wire [63:0] _T_1179; // @[Mux.scala 19:72:Sodor3Stage.fir@2622.4]
  wire [63:0] _GEN_407; // @[Mux.scala 19:72:Sodor3Stage.fir@2623.4]
  wire [63:0] _T_1180; // @[Mux.scala 19:72:Sodor3Stage.fir@2623.4]
  wire [63:0] _GEN_408; // @[Mux.scala 19:72:Sodor3Stage.fir@2624.4]
  wire [63:0] _T_1181; // @[Mux.scala 19:72:Sodor3Stage.fir@2624.4]
  wire [63:0] _GEN_409; // @[Mux.scala 19:72:Sodor3Stage.fir@2625.4]
  wire [63:0] _T_1182; // @[Mux.scala 19:72:Sodor3Stage.fir@2625.4]
  wire [63:0] _GEN_410; // @[Mux.scala 19:72:Sodor3Stage.fir@2626.4]
  wire [63:0] _T_1183; // @[Mux.scala 19:72:Sodor3Stage.fir@2626.4]
  wire [63:0] _GEN_411; // @[Mux.scala 19:72:Sodor3Stage.fir@2627.4]
  wire [63:0] _T_1184; // @[Mux.scala 19:72:Sodor3Stage.fir@2627.4]
  wire [63:0] _GEN_412; // @[Mux.scala 19:72:Sodor3Stage.fir@2628.4]
  wire [63:0] _T_1185; // @[Mux.scala 19:72:Sodor3Stage.fir@2628.4]
  wire [63:0] _GEN_413; // @[Mux.scala 19:72:Sodor3Stage.fir@2629.4]
  wire [63:0] _T_1186; // @[Mux.scala 19:72:Sodor3Stage.fir@2629.4]
  wire [63:0] _GEN_414; // @[Mux.scala 19:72:Sodor3Stage.fir@2630.4]
  wire [63:0] _T_1187; // @[Mux.scala 19:72:Sodor3Stage.fir@2630.4]
  wire [63:0] _GEN_415; // @[Mux.scala 19:72:Sodor3Stage.fir@2631.4]
  wire [63:0] _T_1188; // @[Mux.scala 19:72:Sodor3Stage.fir@2631.4]
  wire [63:0] _GEN_416; // @[Mux.scala 19:72:Sodor3Stage.fir@2632.4]
  wire [63:0] _T_1189; // @[Mux.scala 19:72:Sodor3Stage.fir@2632.4]
  wire [63:0] _GEN_417; // @[Mux.scala 19:72:Sodor3Stage.fir@2633.4]
  wire [63:0] _T_1190; // @[Mux.scala 19:72:Sodor3Stage.fir@2633.4]
  wire [63:0] _GEN_418; // @[Mux.scala 19:72:Sodor3Stage.fir@2634.4]
  wire [63:0] _T_1191; // @[Mux.scala 19:72:Sodor3Stage.fir@2634.4]
  wire [63:0] _GEN_419; // @[Mux.scala 19:72:Sodor3Stage.fir@2635.4]
  wire [63:0] _T_1192; // @[Mux.scala 19:72:Sodor3Stage.fir@2635.4]
  wire [63:0] _GEN_420; // @[Mux.scala 19:72:Sodor3Stage.fir@2636.4]
  wire [63:0] _T_1193; // @[Mux.scala 19:72:Sodor3Stage.fir@2636.4]
  wire [63:0] _GEN_421; // @[Mux.scala 19:72:Sodor3Stage.fir@2637.4]
  wire [63:0] _T_1194; // @[Mux.scala 19:72:Sodor3Stage.fir@2637.4]
  wire [63:0] _GEN_422; // @[Mux.scala 19:72:Sodor3Stage.fir@2638.4]
  wire [63:0] _T_1195; // @[Mux.scala 19:72:Sodor3Stage.fir@2638.4]
  wire [63:0] _GEN_423; // @[Mux.scala 19:72:Sodor3Stage.fir@2639.4]
  wire [63:0] _T_1196; // @[Mux.scala 19:72:Sodor3Stage.fir@2639.4]
  wire [63:0] _GEN_424; // @[Mux.scala 19:72:Sodor3Stage.fir@2640.4]
  wire [63:0] _T_1197; // @[Mux.scala 19:72:Sodor3Stage.fir@2640.4]
  wire [63:0] _GEN_425; // @[Mux.scala 19:72:Sodor3Stage.fir@2641.4]
  wire [63:0] _T_1198; // @[Mux.scala 19:72:Sodor3Stage.fir@2641.4]
  wire [63:0] _GEN_426; // @[Mux.scala 19:72:Sodor3Stage.fir@2642.4]
  wire [63:0] _T_1199; // @[Mux.scala 19:72:Sodor3Stage.fir@2642.4]
  wire [63:0] _GEN_427; // @[Mux.scala 19:72:Sodor3Stage.fir@2643.4]
  wire [63:0] _T_1200; // @[Mux.scala 19:72:Sodor3Stage.fir@2643.4]
  wire [63:0] _GEN_428; // @[Mux.scala 19:72:Sodor3Stage.fir@2644.4]
  wire [63:0] _T_1201; // @[Mux.scala 19:72:Sodor3Stage.fir@2644.4]
  wire [63:0] _GEN_429; // @[Mux.scala 19:72:Sodor3Stage.fir@2645.4]
  wire [63:0] _T_1202; // @[Mux.scala 19:72:Sodor3Stage.fir@2645.4]
  wire [63:0] _GEN_430; // @[Mux.scala 19:72:Sodor3Stage.fir@2646.4]
  wire [63:0] _T_1203; // @[Mux.scala 19:72:Sodor3Stage.fir@2646.4]
  wire [63:0] _GEN_431; // @[Mux.scala 19:72:Sodor3Stage.fir@2647.4]
  wire [63:0] _T_1204; // @[Mux.scala 19:72:Sodor3Stage.fir@2647.4]
  wire [63:0] _GEN_432; // @[Mux.scala 19:72:Sodor3Stage.fir@2648.4]
  wire [63:0] _T_1205; // @[Mux.scala 19:72:Sodor3Stage.fir@2648.4]
  wire [63:0] _GEN_433; // @[Mux.scala 19:72:Sodor3Stage.fir@2649.4]
  wire [63:0] _T_1206; // @[Mux.scala 19:72:Sodor3Stage.fir@2649.4]
  wire [63:0] _GEN_434; // @[Mux.scala 19:72:Sodor3Stage.fir@2650.4]
  wire [63:0] _T_1207; // @[Mux.scala 19:72:Sodor3Stage.fir@2650.4]
  wire [63:0] _GEN_435; // @[Mux.scala 19:72:Sodor3Stage.fir@2651.4]
  wire [63:0] _T_1208; // @[Mux.scala 19:72:Sodor3Stage.fir@2651.4]
  wire [63:0] _GEN_436; // @[Mux.scala 19:72:Sodor3Stage.fir@2652.4]
  wire [63:0] _T_1209; // @[Mux.scala 19:72:Sodor3Stage.fir@2652.4]
  wire [63:0] _GEN_437; // @[Mux.scala 19:72:Sodor3Stage.fir@2653.4]
  wire [63:0] _T_1210; // @[Mux.scala 19:72:Sodor3Stage.fir@2653.4]
  wire [63:0] _GEN_438; // @[Mux.scala 19:72:Sodor3Stage.fir@2654.4]
  wire [63:0] _T_1211; // @[Mux.scala 19:72:Sodor3Stage.fir@2654.4]
  wire [63:0] _GEN_439; // @[Mux.scala 19:72:Sodor3Stage.fir@2655.4]
  wire [63:0] _T_1212; // @[Mux.scala 19:72:Sodor3Stage.fir@2655.4]
  wire [63:0] _GEN_440; // @[Mux.scala 19:72:Sodor3Stage.fir@2656.4]
  wire [63:0] _T_1213; // @[Mux.scala 19:72:Sodor3Stage.fir@2656.4]
  wire [63:0] _GEN_441; // @[Mux.scala 19:72:Sodor3Stage.fir@2657.4]
  wire [63:0] _T_1214; // @[Mux.scala 19:72:Sodor3Stage.fir@2657.4]
  wire [63:0] _GEN_442; // @[Mux.scala 19:72:Sodor3Stage.fir@2658.4]
  wire [63:0] _T_1215; // @[Mux.scala 19:72:Sodor3Stage.fir@2658.4]
  wire [63:0] _GEN_443; // @[Mux.scala 19:72:Sodor3Stage.fir@2659.4]
  wire [63:0] _T_1216; // @[Mux.scala 19:72:Sodor3Stage.fir@2659.4]
  wire [63:0] _GEN_444; // @[Mux.scala 19:72:Sodor3Stage.fir@2660.4]
  wire [63:0] _T_1217; // @[Mux.scala 19:72:Sodor3Stage.fir@2660.4]
  wire [63:0] _GEN_445; // @[Mux.scala 19:72:Sodor3Stage.fir@2661.4]
  wire [63:0] _T_1218; // @[Mux.scala 19:72:Sodor3Stage.fir@2661.4]
  wire [63:0] _GEN_446; // @[Mux.scala 19:72:Sodor3Stage.fir@2662.4]
  wire [63:0] _T_1219; // @[Mux.scala 19:72:Sodor3Stage.fir@2662.4]
  wire [63:0] _GEN_447; // @[Mux.scala 19:72:Sodor3Stage.fir@2663.4]
  wire [63:0] _T_1220; // @[Mux.scala 19:72:Sodor3Stage.fir@2663.4]
  wire [63:0] _GEN_448; // @[Mux.scala 19:72:Sodor3Stage.fir@2664.4]
  wire [63:0] _T_1221; // @[Mux.scala 19:72:Sodor3Stage.fir@2664.4]
  wire [63:0] _GEN_449; // @[Mux.scala 19:72:Sodor3Stage.fir@2665.4]
  wire [63:0] _T_1222; // @[Mux.scala 19:72:Sodor3Stage.fir@2665.4]
  wire [63:0] _GEN_450; // @[Mux.scala 19:72:Sodor3Stage.fir@2666.4]
  wire [63:0] _T_1223; // @[Mux.scala 19:72:Sodor3Stage.fir@2666.4]
  wire [63:0] _GEN_451; // @[Mux.scala 19:72:Sodor3Stage.fir@2667.4]
  wire [63:0] _T_1224; // @[Mux.scala 19:72:Sodor3Stage.fir@2667.4]
  wire [63:0] _GEN_452; // @[Mux.scala 19:72:Sodor3Stage.fir@2668.4]
  wire [63:0] _T_1225; // @[Mux.scala 19:72:Sodor3Stage.fir@2668.4]
  wire [63:0] _GEN_453; // @[Mux.scala 19:72:Sodor3Stage.fir@2669.4]
  wire [63:0] _T_1226; // @[Mux.scala 19:72:Sodor3Stage.fir@2669.4]
  wire [63:0] _GEN_454; // @[Mux.scala 19:72:Sodor3Stage.fir@2670.4]
  wire [63:0] _T_1227; // @[Mux.scala 19:72:Sodor3Stage.fir@2670.4]
  wire [63:0] _GEN_455; // @[Mux.scala 19:72:Sodor3Stage.fir@2671.4]
  wire [63:0] _T_1228; // @[Mux.scala 19:72:Sodor3Stage.fir@2671.4]
  wire [63:0] _GEN_456; // @[Mux.scala 19:72:Sodor3Stage.fir@2672.4]
  wire [63:0] _T_1229; // @[Mux.scala 19:72:Sodor3Stage.fir@2672.4]
  wire [63:0] _GEN_457; // @[Mux.scala 19:72:Sodor3Stage.fir@2673.4]
  wire [63:0] _T_1230; // @[Mux.scala 19:72:Sodor3Stage.fir@2673.4]
  wire [63:0] _GEN_458; // @[Mux.scala 19:72:Sodor3Stage.fir@2674.4]
  wire [63:0] _T_1231; // @[Mux.scala 19:72:Sodor3Stage.fir@2674.4]
  wire [63:0] _GEN_459; // @[Mux.scala 19:72:Sodor3Stage.fir@2675.4]
  wire [63:0] _T_1232; // @[Mux.scala 19:72:Sodor3Stage.fir@2675.4]
  wire [63:0] _GEN_460; // @[Mux.scala 19:72:Sodor3Stage.fir@2676.4]
  wire [63:0] _T_1233; // @[Mux.scala 19:72:Sodor3Stage.fir@2676.4]
  wire [63:0] _GEN_461; // @[Mux.scala 19:72:Sodor3Stage.fir@2677.4]
  wire [63:0] _T_1234; // @[Mux.scala 19:72:Sodor3Stage.fir@2677.4]
  wire [63:0] _GEN_462; // @[Mux.scala 19:72:Sodor3Stage.fir@2678.4]
  wire [63:0] _T_1235; // @[Mux.scala 19:72:Sodor3Stage.fir@2678.4]
  wire [63:0] _GEN_463; // @[Mux.scala 19:72:Sodor3Stage.fir@2679.4]
  wire [63:0] _T_1236; // @[Mux.scala 19:72:Sodor3Stage.fir@2679.4]
  wire [63:0] _GEN_464; // @[Mux.scala 19:72:Sodor3Stage.fir@2680.4]
  wire [63:0] _T_1237; // @[Mux.scala 19:72:Sodor3Stage.fir@2680.4]
  wire [63:0] _GEN_465; // @[Mux.scala 19:72:Sodor3Stage.fir@2681.4]
  wire [63:0] _T_1238; // @[Mux.scala 19:72:Sodor3Stage.fir@2681.4]
  wire [63:0] _GEN_466; // @[Mux.scala 19:72:Sodor3Stage.fir@2682.4]
  wire [63:0] _T_1239; // @[Mux.scala 19:72:Sodor3Stage.fir@2682.4]
  wire [63:0] _GEN_467; // @[Mux.scala 19:72:Sodor3Stage.fir@2683.4]
  wire [63:0] _T_1240; // @[Mux.scala 19:72:Sodor3Stage.fir@2683.4]
  wire [63:0] _GEN_468; // @[Mux.scala 19:72:Sodor3Stage.fir@2684.4]
  wire [63:0] _T_1241; // @[Mux.scala 19:72:Sodor3Stage.fir@2684.4]
  wire  _T_1252; // @[csr.scala 334:43:Sodor3Stage.fir@2697.8]
  wire  _T_1262; // @[csr.scala 334:43:Sodor3Stage.fir@2717.8]
  wire [34:0] _T_1270; // @[:Sodor3Stage.fir@2730.8]
  wire  _T_1274; // @[csr.scala 341:47:Sodor3Stage.fir@2738.8]
  wire  _T_1278; // @[csr.scala 341:47:Sodor3Stage.fir@2746.8]
  wire [15:0] _T_1298; // @[:Sodor3Stage.fir@2783.8]
  wire  _T_1302; // @[csr.scala 346:39:Sodor3Stage.fir@2791.8]
  wire  _T_1306; // @[csr.scala 346:39:Sodor3Stage.fir@2799.8]
  wire [7:0] _T_1336; // @[csr.scala 386:47:Sodor3Stage.fir@2859.8]
  wire [31:0] _T_1337; // @[csr.scala 386:72:Sodor3Stage.fir@2860.8]
  wire [39:0] _T_1338; // @[Cat.scala 30:58:Sodor3Stage.fir@2861.8]
  wire [40:0] _GEN_24; // @[csr.scala 386:29:Sodor3Stage.fir@2858.6]
  wire [7:0] _T_1339; // @[csr.scala 387:45:Sodor3Stage.fir@2865.8]
  wire [39:0] _T_1340; // @[Cat.scala 30:58:Sodor3Stage.fir@2866.8]
  wire [40:0] _GEN_25; // @[csr.scala 387:29:Sodor3Stage.fir@2864.6]
  wire [31:0] _T_1342; // @[csr.scala 386:72:Sodor3Stage.fir@2871.8]
  wire [39:0] _T_1343; // @[Cat.scala 30:58:Sodor3Stage.fir@2872.8]
  wire [40:0] _GEN_26; // @[csr.scala 386:29:Sodor3Stage.fir@2869.6]
  wire [7:0] _T_1344; // @[csr.scala 387:45:Sodor3Stage.fir@2876.8]
  wire [39:0] _T_1345; // @[Cat.scala 30:58:Sodor3Stage.fir@2877.8]
  wire [40:0] _GEN_27; // @[csr.scala 387:29:Sodor3Stage.fir@2875.6]
  wire [31:0] _T_1347; // @[csr.scala 386:72:Sodor3Stage.fir@2882.8]
  wire [39:0] _T_1348; // @[Cat.scala 30:58:Sodor3Stage.fir@2883.8]
  wire [40:0] _GEN_28; // @[csr.scala 386:29:Sodor3Stage.fir@2880.6]
  wire [7:0] _T_1349; // @[csr.scala 387:45:Sodor3Stage.fir@2887.8]
  wire [39:0] _T_1350; // @[Cat.scala 30:58:Sodor3Stage.fir@2888.8]
  wire [40:0] _GEN_29; // @[csr.scala 387:29:Sodor3Stage.fir@2886.6]
  wire [31:0] _T_1352; // @[csr.scala 386:72:Sodor3Stage.fir@2893.8]
  wire [39:0] _T_1353; // @[Cat.scala 30:58:Sodor3Stage.fir@2894.8]
  wire [40:0] _GEN_30; // @[csr.scala 386:29:Sodor3Stage.fir@2891.6]
  wire [7:0] _T_1354; // @[csr.scala 387:45:Sodor3Stage.fir@2898.8]
  wire [39:0] _T_1355; // @[Cat.scala 30:58:Sodor3Stage.fir@2899.8]
  wire [40:0] _GEN_31; // @[csr.scala 387:29:Sodor3Stage.fir@2897.6]
  wire [31:0] _T_1357; // @[csr.scala 386:72:Sodor3Stage.fir@2904.8]
  wire [39:0] _T_1358; // @[Cat.scala 30:58:Sodor3Stage.fir@2905.8]
  wire [40:0] _GEN_32; // @[csr.scala 386:29:Sodor3Stage.fir@2902.6]
  wire [7:0] _T_1359; // @[csr.scala 387:45:Sodor3Stage.fir@2909.8]
  wire [39:0] _T_1360; // @[Cat.scala 30:58:Sodor3Stage.fir@2910.8]
  wire [40:0] _GEN_33; // @[csr.scala 387:29:Sodor3Stage.fir@2908.6]
  wire [31:0] _T_1362; // @[csr.scala 386:72:Sodor3Stage.fir@2915.8]
  wire [39:0] _T_1363; // @[Cat.scala 30:58:Sodor3Stage.fir@2916.8]
  wire [40:0] _GEN_34; // @[csr.scala 386:29:Sodor3Stage.fir@2913.6]
  wire [7:0] _T_1364; // @[csr.scala 387:45:Sodor3Stage.fir@2920.8]
  wire [39:0] _T_1365; // @[Cat.scala 30:58:Sodor3Stage.fir@2921.8]
  wire [40:0] _GEN_35; // @[csr.scala 387:29:Sodor3Stage.fir@2919.6]
  wire [31:0] _T_1367; // @[csr.scala 386:72:Sodor3Stage.fir@2926.8]
  wire [39:0] _T_1368; // @[Cat.scala 30:58:Sodor3Stage.fir@2927.8]
  wire [40:0] _GEN_36; // @[csr.scala 386:29:Sodor3Stage.fir@2924.6]
  wire [7:0] _T_1369; // @[csr.scala 387:45:Sodor3Stage.fir@2931.8]
  wire [39:0] _T_1370; // @[Cat.scala 30:58:Sodor3Stage.fir@2932.8]
  wire [40:0] _GEN_37; // @[csr.scala 387:29:Sodor3Stage.fir@2930.6]
  wire [31:0] _T_1372; // @[csr.scala 386:72:Sodor3Stage.fir@2937.8]
  wire [39:0] _T_1373; // @[Cat.scala 30:58:Sodor3Stage.fir@2938.8]
  wire [40:0] _GEN_38; // @[csr.scala 386:29:Sodor3Stage.fir@2935.6]
  wire [7:0] _T_1374; // @[csr.scala 387:45:Sodor3Stage.fir@2942.8]
  wire [39:0] _T_1375; // @[Cat.scala 30:58:Sodor3Stage.fir@2943.8]
  wire [40:0] _GEN_39; // @[csr.scala 387:29:Sodor3Stage.fir@2941.6]
  wire [31:0] _T_1377; // @[csr.scala 386:72:Sodor3Stage.fir@2948.8]
  wire [39:0] _T_1378; // @[Cat.scala 30:58:Sodor3Stage.fir@2949.8]
  wire [40:0] _GEN_40; // @[csr.scala 386:29:Sodor3Stage.fir@2946.6]
  wire [7:0] _T_1379; // @[csr.scala 387:45:Sodor3Stage.fir@2953.8]
  wire [39:0] _T_1380; // @[Cat.scala 30:58:Sodor3Stage.fir@2954.8]
  wire [40:0] _GEN_41; // @[csr.scala 387:29:Sodor3Stage.fir@2952.6]
  wire [31:0] _T_1382; // @[csr.scala 386:72:Sodor3Stage.fir@2959.8]
  wire [39:0] _T_1383; // @[Cat.scala 30:58:Sodor3Stage.fir@2960.8]
  wire [40:0] _GEN_42; // @[csr.scala 386:29:Sodor3Stage.fir@2957.6]
  wire [7:0] _T_1384; // @[csr.scala 387:45:Sodor3Stage.fir@2964.8]
  wire [39:0] _T_1385; // @[Cat.scala 30:58:Sodor3Stage.fir@2965.8]
  wire [40:0] _GEN_43; // @[csr.scala 387:29:Sodor3Stage.fir@2963.6]
  wire [31:0] _T_1387; // @[csr.scala 386:72:Sodor3Stage.fir@2970.8]
  wire [39:0] _T_1388; // @[Cat.scala 30:58:Sodor3Stage.fir@2971.8]
  wire [40:0] _GEN_44; // @[csr.scala 386:29:Sodor3Stage.fir@2968.6]
  wire [7:0] _T_1389; // @[csr.scala 387:45:Sodor3Stage.fir@2975.8]
  wire [39:0] _T_1390; // @[Cat.scala 30:58:Sodor3Stage.fir@2976.8]
  wire [40:0] _GEN_45; // @[csr.scala 387:29:Sodor3Stage.fir@2974.6]
  wire [31:0] _T_1392; // @[csr.scala 386:72:Sodor3Stage.fir@2981.8]
  wire [39:0] _T_1393; // @[Cat.scala 30:58:Sodor3Stage.fir@2982.8]
  wire [40:0] _GEN_46; // @[csr.scala 386:29:Sodor3Stage.fir@2979.6]
  wire [7:0] _T_1394; // @[csr.scala 387:45:Sodor3Stage.fir@2986.8]
  wire [39:0] _T_1395; // @[Cat.scala 30:58:Sodor3Stage.fir@2987.8]
  wire [40:0] _GEN_47; // @[csr.scala 387:29:Sodor3Stage.fir@2985.6]
  wire [31:0] _T_1397; // @[csr.scala 386:72:Sodor3Stage.fir@2992.8]
  wire [39:0] _T_1398; // @[Cat.scala 30:58:Sodor3Stage.fir@2993.8]
  wire [40:0] _GEN_48; // @[csr.scala 386:29:Sodor3Stage.fir@2990.6]
  wire [7:0] _T_1399; // @[csr.scala 387:45:Sodor3Stage.fir@2997.8]
  wire [39:0] _T_1400; // @[Cat.scala 30:58:Sodor3Stage.fir@2998.8]
  wire [40:0] _GEN_49; // @[csr.scala 387:29:Sodor3Stage.fir@2996.6]
  wire [31:0] _T_1402; // @[csr.scala 386:72:Sodor3Stage.fir@3003.8]
  wire [39:0] _T_1403; // @[Cat.scala 30:58:Sodor3Stage.fir@3004.8]
  wire [40:0] _GEN_50; // @[csr.scala 386:29:Sodor3Stage.fir@3001.6]
  wire [7:0] _T_1404; // @[csr.scala 387:45:Sodor3Stage.fir@3008.8]
  wire [39:0] _T_1405; // @[Cat.scala 30:58:Sodor3Stage.fir@3009.8]
  wire [40:0] _GEN_51; // @[csr.scala 387:29:Sodor3Stage.fir@3007.6]
  wire [31:0] _T_1407; // @[csr.scala 386:72:Sodor3Stage.fir@3014.8]
  wire [39:0] _T_1408; // @[Cat.scala 30:58:Sodor3Stage.fir@3015.8]
  wire [40:0] _GEN_52; // @[csr.scala 386:29:Sodor3Stage.fir@3012.6]
  wire [7:0] _T_1409; // @[csr.scala 387:45:Sodor3Stage.fir@3019.8]
  wire [39:0] _T_1410; // @[Cat.scala 30:58:Sodor3Stage.fir@3020.8]
  wire [40:0] _GEN_53; // @[csr.scala 387:29:Sodor3Stage.fir@3018.6]
  wire [31:0] _T_1412; // @[csr.scala 386:72:Sodor3Stage.fir@3025.8]
  wire [39:0] _T_1413; // @[Cat.scala 30:58:Sodor3Stage.fir@3026.8]
  wire [40:0] _GEN_54; // @[csr.scala 386:29:Sodor3Stage.fir@3023.6]
  wire [7:0] _T_1414; // @[csr.scala 387:45:Sodor3Stage.fir@3030.8]
  wire [39:0] _T_1415; // @[Cat.scala 30:58:Sodor3Stage.fir@3031.8]
  wire [40:0] _GEN_55; // @[csr.scala 387:29:Sodor3Stage.fir@3029.6]
  wire [31:0] _T_1417; // @[csr.scala 386:72:Sodor3Stage.fir@3036.8]
  wire [39:0] _T_1418; // @[Cat.scala 30:58:Sodor3Stage.fir@3037.8]
  wire [40:0] _GEN_56; // @[csr.scala 386:29:Sodor3Stage.fir@3034.6]
  wire [7:0] _T_1419; // @[csr.scala 387:45:Sodor3Stage.fir@3041.8]
  wire [39:0] _T_1420; // @[Cat.scala 30:58:Sodor3Stage.fir@3042.8]
  wire [40:0] _GEN_57; // @[csr.scala 387:29:Sodor3Stage.fir@3040.6]
  wire [31:0] _T_1422; // @[csr.scala 386:72:Sodor3Stage.fir@3047.8]
  wire [39:0] _T_1423; // @[Cat.scala 30:58:Sodor3Stage.fir@3048.8]
  wire [40:0] _GEN_58; // @[csr.scala 386:29:Sodor3Stage.fir@3045.6]
  wire [7:0] _T_1424; // @[csr.scala 387:45:Sodor3Stage.fir@3052.8]
  wire [39:0] _T_1425; // @[Cat.scala 30:58:Sodor3Stage.fir@3053.8]
  wire [40:0] _GEN_59; // @[csr.scala 387:29:Sodor3Stage.fir@3051.6]
  wire [31:0] _T_1427; // @[csr.scala 386:72:Sodor3Stage.fir@3058.8]
  wire [39:0] _T_1428; // @[Cat.scala 30:58:Sodor3Stage.fir@3059.8]
  wire [40:0] _GEN_60; // @[csr.scala 386:29:Sodor3Stage.fir@3056.6]
  wire [7:0] _T_1429; // @[csr.scala 387:45:Sodor3Stage.fir@3063.8]
  wire [39:0] _T_1430; // @[Cat.scala 30:58:Sodor3Stage.fir@3064.8]
  wire [40:0] _GEN_61; // @[csr.scala 387:29:Sodor3Stage.fir@3062.6]
  wire [31:0] _T_1432; // @[csr.scala 386:72:Sodor3Stage.fir@3069.8]
  wire [39:0] _T_1433; // @[Cat.scala 30:58:Sodor3Stage.fir@3070.8]
  wire [40:0] _GEN_62; // @[csr.scala 386:29:Sodor3Stage.fir@3067.6]
  wire [7:0] _T_1434; // @[csr.scala 387:45:Sodor3Stage.fir@3074.8]
  wire [39:0] _T_1435; // @[Cat.scala 30:58:Sodor3Stage.fir@3075.8]
  wire [40:0] _GEN_63; // @[csr.scala 387:29:Sodor3Stage.fir@3073.6]
  wire [31:0] _T_1437; // @[csr.scala 386:72:Sodor3Stage.fir@3080.8]
  wire [39:0] _T_1438; // @[Cat.scala 30:58:Sodor3Stage.fir@3081.8]
  wire [40:0] _GEN_64; // @[csr.scala 386:29:Sodor3Stage.fir@3078.6]
  wire [7:0] _T_1439; // @[csr.scala 387:45:Sodor3Stage.fir@3085.8]
  wire [39:0] _T_1440; // @[Cat.scala 30:58:Sodor3Stage.fir@3086.8]
  wire [40:0] _GEN_65; // @[csr.scala 387:29:Sodor3Stage.fir@3084.6]
  wire [31:0] _T_1442; // @[csr.scala 386:72:Sodor3Stage.fir@3091.8]
  wire [39:0] _T_1443; // @[Cat.scala 30:58:Sodor3Stage.fir@3092.8]
  wire [40:0] _GEN_66; // @[csr.scala 386:29:Sodor3Stage.fir@3089.6]
  wire [7:0] _T_1444; // @[csr.scala 387:45:Sodor3Stage.fir@3096.8]
  wire [39:0] _T_1445; // @[Cat.scala 30:58:Sodor3Stage.fir@3097.8]
  wire [40:0] _GEN_67; // @[csr.scala 387:29:Sodor3Stage.fir@3095.6]
  wire [31:0] _T_1447; // @[csr.scala 386:72:Sodor3Stage.fir@3102.8]
  wire [39:0] _T_1448; // @[Cat.scala 30:58:Sodor3Stage.fir@3103.8]
  wire [40:0] _GEN_68; // @[csr.scala 386:29:Sodor3Stage.fir@3100.6]
  wire [7:0] _T_1449; // @[csr.scala 387:45:Sodor3Stage.fir@3107.8]
  wire [39:0] _T_1450; // @[Cat.scala 30:58:Sodor3Stage.fir@3108.8]
  wire [40:0] _GEN_69; // @[csr.scala 387:29:Sodor3Stage.fir@3106.6]
  wire [31:0] _T_1452; // @[csr.scala 386:72:Sodor3Stage.fir@3113.8]
  wire [39:0] _T_1453; // @[Cat.scala 30:58:Sodor3Stage.fir@3114.8]
  wire [40:0] _GEN_70; // @[csr.scala 386:29:Sodor3Stage.fir@3111.6]
  wire [7:0] _T_1454; // @[csr.scala 387:45:Sodor3Stage.fir@3118.8]
  wire [39:0] _T_1455; // @[Cat.scala 30:58:Sodor3Stage.fir@3119.8]
  wire [40:0] _GEN_71; // @[csr.scala 387:29:Sodor3Stage.fir@3117.6]
  wire [31:0] _T_1457; // @[csr.scala 386:72:Sodor3Stage.fir@3124.8]
  wire [39:0] _T_1458; // @[Cat.scala 30:58:Sodor3Stage.fir@3125.8]
  wire [40:0] _GEN_72; // @[csr.scala 386:29:Sodor3Stage.fir@3122.6]
  wire [7:0] _T_1459; // @[csr.scala 387:45:Sodor3Stage.fir@3129.8]
  wire [39:0] _T_1460; // @[Cat.scala 30:58:Sodor3Stage.fir@3130.8]
  wire [40:0] _GEN_73; // @[csr.scala 387:29:Sodor3Stage.fir@3128.6]
  wire [31:0] _T_1462; // @[csr.scala 386:72:Sodor3Stage.fir@3135.8]
  wire [39:0] _T_1463; // @[Cat.scala 30:58:Sodor3Stage.fir@3136.8]
  wire [40:0] _GEN_74; // @[csr.scala 386:29:Sodor3Stage.fir@3133.6]
  wire [7:0] _T_1464; // @[csr.scala 387:45:Sodor3Stage.fir@3140.8]
  wire [39:0] _T_1465; // @[Cat.scala 30:58:Sodor3Stage.fir@3141.8]
  wire [40:0] _GEN_75; // @[csr.scala 387:29:Sodor3Stage.fir@3139.6]
  wire [31:0] _T_1467; // @[csr.scala 386:72:Sodor3Stage.fir@3146.8]
  wire [39:0] _T_1468; // @[Cat.scala 30:58:Sodor3Stage.fir@3147.8]
  wire [40:0] _GEN_76; // @[csr.scala 386:29:Sodor3Stage.fir@3144.6]
  wire [7:0] _T_1469; // @[csr.scala 387:45:Sodor3Stage.fir@3151.8]
  wire [39:0] _T_1470; // @[Cat.scala 30:58:Sodor3Stage.fir@3152.8]
  wire [40:0] _GEN_77; // @[csr.scala 387:29:Sodor3Stage.fir@3150.6]
  wire [31:0] _T_1472; // @[csr.scala 386:72:Sodor3Stage.fir@3157.8]
  wire [39:0] _T_1473; // @[Cat.scala 30:58:Sodor3Stage.fir@3158.8]
  wire [40:0] _GEN_78; // @[csr.scala 386:29:Sodor3Stage.fir@3155.6]
  wire [7:0] _T_1474; // @[csr.scala 387:45:Sodor3Stage.fir@3162.8]
  wire [39:0] _T_1475; // @[Cat.scala 30:58:Sodor3Stage.fir@3163.8]
  wire [40:0] _GEN_79; // @[csr.scala 387:29:Sodor3Stage.fir@3161.6]
  wire [31:0] _T_1477; // @[csr.scala 386:72:Sodor3Stage.fir@3168.8]
  wire [39:0] _T_1478; // @[Cat.scala 30:58:Sodor3Stage.fir@3169.8]
  wire [40:0] _GEN_80; // @[csr.scala 386:29:Sodor3Stage.fir@3166.6]
  wire [7:0] _T_1479; // @[csr.scala 387:45:Sodor3Stage.fir@3173.8]
  wire [39:0] _T_1480; // @[Cat.scala 30:58:Sodor3Stage.fir@3174.8]
  wire [40:0] _GEN_81; // @[csr.scala 387:29:Sodor3Stage.fir@3172.6]
  wire [31:0] _T_1482; // @[csr.scala 386:72:Sodor3Stage.fir@3179.8]
  wire [39:0] _T_1483; // @[Cat.scala 30:58:Sodor3Stage.fir@3180.8]
  wire [40:0] _GEN_82; // @[csr.scala 386:29:Sodor3Stage.fir@3177.6]
  wire [7:0] _T_1484; // @[csr.scala 387:45:Sodor3Stage.fir@3184.8]
  wire [39:0] _T_1485; // @[Cat.scala 30:58:Sodor3Stage.fir@3185.8]
  wire [40:0] _GEN_83; // @[csr.scala 387:29:Sodor3Stage.fir@3183.6]
  wire [31:0] _T_1487; // @[csr.scala 386:72:Sodor3Stage.fir@3190.8]
  wire [39:0] _T_1488; // @[Cat.scala 30:58:Sodor3Stage.fir@3191.8]
  wire [40:0] _GEN_84; // @[csr.scala 386:29:Sodor3Stage.fir@3188.6]
  wire [7:0] _T_1489; // @[csr.scala 387:45:Sodor3Stage.fir@3195.8]
  wire [39:0] _T_1490; // @[Cat.scala 30:58:Sodor3Stage.fir@3196.8]
  wire [40:0] _GEN_85; // @[csr.scala 387:29:Sodor3Stage.fir@3194.6]
  wire [31:0] _T_1492; // @[csr.scala 386:72:Sodor3Stage.fir@3201.8]
  wire [39:0] _T_1493; // @[Cat.scala 30:58:Sodor3Stage.fir@3202.8]
  wire [40:0] _GEN_86; // @[csr.scala 386:29:Sodor3Stage.fir@3199.6]
  wire [7:0] _T_1494; // @[csr.scala 387:45:Sodor3Stage.fir@3206.8]
  wire [39:0] _T_1495; // @[Cat.scala 30:58:Sodor3Stage.fir@3207.8]
  wire [40:0] _GEN_87; // @[csr.scala 387:29:Sodor3Stage.fir@3205.6]
  wire [31:0] _T_1497; // @[csr.scala 386:72:Sodor3Stage.fir@3212.8]
  wire [63:0] _T_1498; // @[Cat.scala 30:58:Sodor3Stage.fir@3213.8]
  wire [57:0] _T_1499; // @[util.scala 135:28:Sodor3Stage.fir@3215.8]
  wire [63:0] _GEN_88; // @[csr.scala 386:29:Sodor3Stage.fir@3210.6]
  wire [31:0] _T_1500; // @[csr.scala 387:45:Sodor3Stage.fir@3219.8]
  wire [63:0] _T_1501; // @[Cat.scala 30:58:Sodor3Stage.fir@3220.8]
  wire [57:0] _T_1502; // @[util.scala 135:28:Sodor3Stage.fir@3222.8]
  wire [63:0] _GEN_90; // @[csr.scala 387:29:Sodor3Stage.fir@3218.6]
  wire [31:0] _T_1504; // @[csr.scala 386:72:Sodor3Stage.fir@3227.8]
  wire [63:0] _T_1505; // @[Cat.scala 30:58:Sodor3Stage.fir@3228.8]
  wire [57:0] _T_1506; // @[util.scala 135:28:Sodor3Stage.fir@3230.8]
  wire [63:0] _GEN_92; // @[csr.scala 386:29:Sodor3Stage.fir@3225.6]
  wire [31:0] _T_1507; // @[csr.scala 387:45:Sodor3Stage.fir@3234.8]
  wire [63:0] _T_1508; // @[Cat.scala 30:58:Sodor3Stage.fir@3235.8]
  wire [57:0] _T_1509; // @[util.scala 135:28:Sodor3Stage.fir@3237.8]
  wire [63:0] _GEN_94; // @[csr.scala 387:29:Sodor3Stage.fir@3233.6]
  wire [31:0] _T_1512; // @[csr.scala 368:78:Sodor3Stage.fir@3248.8]
  wire [34:0] _GEN_469; // @[csr.scala 368:86:Sodor3Stage.fir@3249.8]
  wire [34:0] _T_1514; // @[csr.scala 368:86:Sodor3Stage.fir@3249.8]
  wire [34:0] _GEN_98; // @[csr.scala 368:40:Sodor3Stage.fir@3246.6]
  wire [31:0] _T_1516; // @[csr.scala 370:62:Sodor3Stage.fir@3256.8]
  wire [40:0] _GEN_110; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_111; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_112; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_113; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_114; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_115; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_116; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_117; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_118; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_119; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_120; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_121; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_122; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_123; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_124; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_125; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_126; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_127; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_128; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_129; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_130; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_131; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_132; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_133; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_134; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_135; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_136; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_137; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_138; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_139; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_140; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [40:0] _GEN_141; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [63:0] _GEN_142; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [63:0] _GEN_144; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  wire [34:0] _GEN_148; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _T_177 = _T_176 + 6'h1; // @[util.scala 115:33:Sodor3Stage.fir@1808.4]
  assign _T_181 = _T_177[6]; // @[util.scala 120:20:Sodor3Stage.fir@1811.4]
  assign _T_183 = _T_180 + 58'h1; // @[util.scala 120:43:Sodor3Stage.fir@1813.6]
  assign _T_184 = _T_183[57:0]; // @[util.scala 120:43:Sodor3Stage.fir@1814.6]
  assign _T_185 = {_T_180,_T_176}; // @[Cat.scala 30:58:Sodor3Stage.fir@1817.4]
  assign _GEN_389 = {{5'd0}, io_retire}; // @[util.scala 115:33:Sodor3Stage.fir@1819.4]
  assign _T_189 = _T_188 + _GEN_389; // @[util.scala 115:33:Sodor3Stage.fir@1819.4]
  assign _T_193 = _T_189[6]; // @[util.scala 120:20:Sodor3Stage.fir@1822.4]
  assign _T_195 = _T_192 + 58'h1; // @[util.scala 120:43:Sodor3Stage.fir@1824.6]
  assign _T_196 = _T_195[57:0]; // @[util.scala 120:43:Sodor3Stage.fir@1825.6]
  assign _T_197 = {_T_192,_T_188}; // @[Cat.scala 30:58:Sodor3Stage.fir@1828.4]
  assign _T_201 = _T_200 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1831.4]
  assign _T_204 = _T_203 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1834.4]
  assign _T_207 = _T_206 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1837.4]
  assign _T_210 = _T_209 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1840.4]
  assign _T_213 = _T_212 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1843.4]
  assign _T_216 = _T_215 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1846.4]
  assign _T_219 = _T_218 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1849.4]
  assign _T_222 = _T_221 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1852.4]
  assign _T_225 = _T_224 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1855.4]
  assign _T_228 = _T_227 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1858.4]
  assign _T_231 = _T_230 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1861.4]
  assign _T_234 = _T_233 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1864.4]
  assign _T_237 = _T_236 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1867.4]
  assign _T_240 = _T_239 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1870.4]
  assign _T_243 = _T_242 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1873.4]
  assign _T_246 = _T_245 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1876.4]
  assign _T_249 = _T_248 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1879.4]
  assign _T_252 = _T_251 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1882.4]
  assign _T_255 = _T_254 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1885.4]
  assign _T_258 = _T_257 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1888.4]
  assign _T_261 = _T_260 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1891.4]
  assign _T_264 = _T_263 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1894.4]
  assign _T_267 = _T_266 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1897.4]
  assign _T_270 = _T_269 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1900.4]
  assign _T_273 = _T_272 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1903.4]
  assign _T_276 = _T_275 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1906.4]
  assign _T_279 = _T_278 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1909.4]
  assign _T_282 = _T_281 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1912.4]
  assign _T_285 = _T_284 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1915.4]
  assign _T_288 = _T_287 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1918.4]
  assign _T_291 = _T_290 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1921.4]
  assign _T_294 = _T_293 + 40'h0; // @[util.scala 115:33:Sodor3Stage.fir@1924.4]
  assign system_insn = io_rw_cmd == 3'h4; // @[csr.scala 196:31:Sodor3Stage.fir@2069.4]
  assign _T_410 = io_rw_cmd != 3'h0; // @[csr.scala 197:27:Sodor3Stage.fir@2070.4]
  assign _T_412 = system_insn == 1'h0; // @[csr.scala 197:39:Sodor3Stage.fir@2071.4]
  assign cpu_ren = _T_410 & _T_412; // @[csr.scala 197:36:Sodor3Stage.fir@2072.4]
  assign _T_413 = {io_status_sie,io_status_uie}; // @[:Sodor3Stage.fir@2073.4]
  assign _T_414 = {io_status_upie,io_status_mie}; // @[:Sodor3Stage.fir@2074.4]
  assign _T_415 = {_T_414,io_status_hie}; // @[:Sodor3Stage.fir@2075.4]
  assign _T_416 = {_T_415,_T_413}; // @[:Sodor3Stage.fir@2076.4]
  assign _T_417 = {io_status_mpie,io_status_hpie}; // @[:Sodor3Stage.fir@2077.4]
  assign _T_418 = {_T_417,io_status_spie}; // @[:Sodor3Stage.fir@2078.4]
  assign _T_419 = {io_status_mpp,io_status_hpp}; // @[:Sodor3Stage.fir@2079.4]
  assign _T_420 = {_T_419,io_status_spp}; // @[:Sodor3Stage.fir@2080.4]
  assign _T_421 = {_T_420,_T_418}; // @[:Sodor3Stage.fir@2081.4]
  assign _T_422 = {_T_421,_T_416}; // @[:Sodor3Stage.fir@2082.4]
  assign _T_423 = {io_status_mprv,io_status_xs}; // @[:Sodor3Stage.fir@2083.4]
  assign _T_424 = {_T_423,io_status_fs}; // @[:Sodor3Stage.fir@2084.4]
  assign _T_425 = {io_status_tvm,io_status_mxr}; // @[:Sodor3Stage.fir@2085.4]
  assign _T_426 = {_T_425,io_status_sum}; // @[:Sodor3Stage.fir@2086.4]
  assign _T_427 = {_T_426,_T_424}; // @[:Sodor3Stage.fir@2087.4]
  assign _T_428 = {io_status_zero1,io_status_tsr}; // @[:Sodor3Stage.fir@2088.4]
  assign _T_429 = {_T_428,io_status_tw}; // @[:Sodor3Stage.fir@2089.4]
  assign _T_430 = {io_status_debug,io_status_prv}; // @[:Sodor3Stage.fir@2090.4]
  assign _T_431 = {_T_430,io_status_sd}; // @[:Sodor3Stage.fir@2091.4]
  assign _T_432 = {_T_431,_T_429}; // @[:Sodor3Stage.fir@2092.4]
  assign _T_433 = {_T_432,_T_427}; // @[:Sodor3Stage.fir@2093.4]
  assign read_mstatus = {_T_433,_T_422}; // @[:Sodor3Stage.fir@2094.4]
  assign _T_441 = {reg_mip_msip,1'h0}; // @[:Sodor3Stage.fir@2096.4]
  assign _T_442 = {_T_441,2'h0}; // @[:Sodor3Stage.fir@2097.4]
  assign _T_444 = {reg_mip_mtip,1'h0}; // @[:Sodor3Stage.fir@2099.4]
  assign _T_445 = {_T_444,2'h0}; // @[:Sodor3Stage.fir@2100.4]
  assign _T_446 = {_T_445,_T_442}; // @[:Sodor3Stage.fir@2101.4]
  assign _T_454 = {8'h0,_T_446}; // @[:Sodor3Stage.fir@2109.4]
  assign _T_456 = {reg_mie_msip,1'h0}; // @[:Sodor3Stage.fir@2111.4]
  assign _T_457 = {_T_456,2'h0}; // @[:Sodor3Stage.fir@2112.4]
  assign _T_459 = {reg_mie_mtip,1'h0}; // @[:Sodor3Stage.fir@2114.4]
  assign _T_460 = {_T_459,2'h0}; // @[:Sodor3Stage.fir@2115.4]
  assign _T_461 = {_T_460,_T_457}; // @[:Sodor3Stage.fir@2116.4]
  assign _T_469 = {8'h0,_T_461}; // @[:Sodor3Stage.fir@2124.4]
  assign _T_470 = {2'h0,reg_dcsr_step}; // @[csr.scala 222:27:Sodor3Stage.fir@2125.4]
  assign _T_471 = {_T_470,2'h3}; // @[csr.scala 222:27:Sodor3Stage.fir@2126.4]
  assign _T_475 = {6'h0,_T_471}; // @[csr.scala 222:27:Sodor3Stage.fir@2130.4]
  assign _T_479 = {12'h0,reg_dcsr_ebreakm}; // @[csr.scala 222:27:Sodor3Stage.fir@2134.4]
  assign _T_481 = {4'h4,_T_479}; // @[csr.scala 222:27:Sodor3Stage.fir@2136.4]
  assign _T_482 = {_T_481,4'h0}; // @[csr.scala 222:27:Sodor3Stage.fir@2137.4]
  assign _T_483 = {_T_482,_T_475}; // @[csr.scala 222:27:Sodor3Stage.fir@2138.4]
  assign _T_487 = io_decode_csr == 12'hb00; // @[csr.scala 259:76:Sodor3Stage.fir@2139.4]
  assign _T_489 = io_decode_csr == 12'hb02; // @[csr.scala 259:76:Sodor3Stage.fir@2140.4]
  assign _T_491 = io_decode_csr == 12'hf13; // @[csr.scala 259:76:Sodor3Stage.fir@2141.4]
  assign _T_497 = io_decode_csr == 12'h301; // @[csr.scala 259:76:Sodor3Stage.fir@2144.4]
  assign _T_499 = io_decode_csr == 12'h300; // @[csr.scala 259:76:Sodor3Stage.fir@2145.4]
  assign _T_501 = io_decode_csr == 12'h305; // @[csr.scala 259:76:Sodor3Stage.fir@2146.4]
  assign _T_503 = io_decode_csr == 12'h344; // @[csr.scala 259:76:Sodor3Stage.fir@2147.4]
  assign _T_505 = io_decode_csr == 12'h304; // @[csr.scala 259:76:Sodor3Stage.fir@2148.4]
  assign _T_507 = io_decode_csr == 12'h340; // @[csr.scala 259:76:Sodor3Stage.fir@2149.4]
  assign _T_509 = io_decode_csr == 12'h341; // @[csr.scala 259:76:Sodor3Stage.fir@2150.4]
  assign _T_511 = io_decode_csr == 12'h343; // @[csr.scala 259:76:Sodor3Stage.fir@2151.4]
  assign _T_513 = io_decode_csr == 12'h342; // @[csr.scala 259:76:Sodor3Stage.fir@2152.4]
  assign _T_517 = io_decode_csr == 12'h7b0; // @[csr.scala 259:76:Sodor3Stage.fir@2154.4]
  assign _T_519 = io_decode_csr == 12'h7b1; // @[csr.scala 259:76:Sodor3Stage.fir@2155.4]
  assign _T_521 = io_decode_csr == 12'h7b2; // @[csr.scala 259:76:Sodor3Stage.fir@2156.4]
  assign _T_523 = io_decode_csr == 12'h302; // @[csr.scala 259:76:Sodor3Stage.fir@2157.4]
  assign _T_525 = io_decode_csr == 12'hb03; // @[csr.scala 259:76:Sodor3Stage.fir@2158.4]
  assign _T_527 = io_decode_csr == 12'hb83; // @[csr.scala 259:76:Sodor3Stage.fir@2159.4]
  assign _T_529 = io_decode_csr == 12'hb04; // @[csr.scala 259:76:Sodor3Stage.fir@2160.4]
  assign _T_531 = io_decode_csr == 12'hb84; // @[csr.scala 259:76:Sodor3Stage.fir@2161.4]
  assign _T_533 = io_decode_csr == 12'hb05; // @[csr.scala 259:76:Sodor3Stage.fir@2162.4]
  assign _T_535 = io_decode_csr == 12'hb85; // @[csr.scala 259:76:Sodor3Stage.fir@2163.4]
  assign _T_537 = io_decode_csr == 12'hb06; // @[csr.scala 259:76:Sodor3Stage.fir@2164.4]
  assign _T_539 = io_decode_csr == 12'hb86; // @[csr.scala 259:76:Sodor3Stage.fir@2165.4]
  assign _T_541 = io_decode_csr == 12'hb07; // @[csr.scala 259:76:Sodor3Stage.fir@2166.4]
  assign _T_543 = io_decode_csr == 12'hb87; // @[csr.scala 259:76:Sodor3Stage.fir@2167.4]
  assign _T_545 = io_decode_csr == 12'hb08; // @[csr.scala 259:76:Sodor3Stage.fir@2168.4]
  assign _T_547 = io_decode_csr == 12'hb88; // @[csr.scala 259:76:Sodor3Stage.fir@2169.4]
  assign _T_549 = io_decode_csr == 12'hb09; // @[csr.scala 259:76:Sodor3Stage.fir@2170.4]
  assign _T_551 = io_decode_csr == 12'hb89; // @[csr.scala 259:76:Sodor3Stage.fir@2171.4]
  assign _T_553 = io_decode_csr == 12'hb0a; // @[csr.scala 259:76:Sodor3Stage.fir@2172.4]
  assign _T_555 = io_decode_csr == 12'hb8a; // @[csr.scala 259:76:Sodor3Stage.fir@2173.4]
  assign _T_557 = io_decode_csr == 12'hb0b; // @[csr.scala 259:76:Sodor3Stage.fir@2174.4]
  assign _T_559 = io_decode_csr == 12'hb8b; // @[csr.scala 259:76:Sodor3Stage.fir@2175.4]
  assign _T_561 = io_decode_csr == 12'hb0c; // @[csr.scala 259:76:Sodor3Stage.fir@2176.4]
  assign _T_563 = io_decode_csr == 12'hb8c; // @[csr.scala 259:76:Sodor3Stage.fir@2177.4]
  assign _T_565 = io_decode_csr == 12'hb0d; // @[csr.scala 259:76:Sodor3Stage.fir@2178.4]
  assign _T_567 = io_decode_csr == 12'hb8d; // @[csr.scala 259:76:Sodor3Stage.fir@2179.4]
  assign _T_569 = io_decode_csr == 12'hb0e; // @[csr.scala 259:76:Sodor3Stage.fir@2180.4]
  assign _T_571 = io_decode_csr == 12'hb8e; // @[csr.scala 259:76:Sodor3Stage.fir@2181.4]
  assign _T_573 = io_decode_csr == 12'hb0f; // @[csr.scala 259:76:Sodor3Stage.fir@2182.4]
  assign _T_575 = io_decode_csr == 12'hb8f; // @[csr.scala 259:76:Sodor3Stage.fir@2183.4]
  assign _T_577 = io_decode_csr == 12'hb10; // @[csr.scala 259:76:Sodor3Stage.fir@2184.4]
  assign _T_579 = io_decode_csr == 12'hb90; // @[csr.scala 259:76:Sodor3Stage.fir@2185.4]
  assign _T_581 = io_decode_csr == 12'hb11; // @[csr.scala 259:76:Sodor3Stage.fir@2186.4]
  assign _T_583 = io_decode_csr == 12'hb91; // @[csr.scala 259:76:Sodor3Stage.fir@2187.4]
  assign _T_585 = io_decode_csr == 12'hb12; // @[csr.scala 259:76:Sodor3Stage.fir@2188.4]
  assign _T_587 = io_decode_csr == 12'hb92; // @[csr.scala 259:76:Sodor3Stage.fir@2189.4]
  assign _T_589 = io_decode_csr == 12'hb13; // @[csr.scala 259:76:Sodor3Stage.fir@2190.4]
  assign _T_591 = io_decode_csr == 12'hb93; // @[csr.scala 259:76:Sodor3Stage.fir@2191.4]
  assign _T_593 = io_decode_csr == 12'hb14; // @[csr.scala 259:76:Sodor3Stage.fir@2192.4]
  assign _T_595 = io_decode_csr == 12'hb94; // @[csr.scala 259:76:Sodor3Stage.fir@2193.4]
  assign _T_597 = io_decode_csr == 12'hb15; // @[csr.scala 259:76:Sodor3Stage.fir@2194.4]
  assign _T_599 = io_decode_csr == 12'hb95; // @[csr.scala 259:76:Sodor3Stage.fir@2195.4]
  assign _T_601 = io_decode_csr == 12'hb16; // @[csr.scala 259:76:Sodor3Stage.fir@2196.4]
  assign _T_603 = io_decode_csr == 12'hb96; // @[csr.scala 259:76:Sodor3Stage.fir@2197.4]
  assign _T_605 = io_decode_csr == 12'hb17; // @[csr.scala 259:76:Sodor3Stage.fir@2198.4]
  assign _T_607 = io_decode_csr == 12'hb97; // @[csr.scala 259:76:Sodor3Stage.fir@2199.4]
  assign _T_609 = io_decode_csr == 12'hb18; // @[csr.scala 259:76:Sodor3Stage.fir@2200.4]
  assign _T_611 = io_decode_csr == 12'hb98; // @[csr.scala 259:76:Sodor3Stage.fir@2201.4]
  assign _T_613 = io_decode_csr == 12'hb19; // @[csr.scala 259:76:Sodor3Stage.fir@2202.4]
  assign _T_615 = io_decode_csr == 12'hb99; // @[csr.scala 259:76:Sodor3Stage.fir@2203.4]
  assign _T_617 = io_decode_csr == 12'hb1a; // @[csr.scala 259:76:Sodor3Stage.fir@2204.4]
  assign _T_619 = io_decode_csr == 12'hb9a; // @[csr.scala 259:76:Sodor3Stage.fir@2205.4]
  assign _T_621 = io_decode_csr == 12'hb1b; // @[csr.scala 259:76:Sodor3Stage.fir@2206.4]
  assign _T_623 = io_decode_csr == 12'hb9b; // @[csr.scala 259:76:Sodor3Stage.fir@2207.4]
  assign _T_625 = io_decode_csr == 12'hb1c; // @[csr.scala 259:76:Sodor3Stage.fir@2208.4]
  assign _T_627 = io_decode_csr == 12'hb9c; // @[csr.scala 259:76:Sodor3Stage.fir@2209.4]
  assign _T_629 = io_decode_csr == 12'hb1d; // @[csr.scala 259:76:Sodor3Stage.fir@2210.4]
  assign _T_631 = io_decode_csr == 12'hb9d; // @[csr.scala 259:76:Sodor3Stage.fir@2211.4]
  assign _T_633 = io_decode_csr == 12'hb1e; // @[csr.scala 259:76:Sodor3Stage.fir@2212.4]
  assign _T_635 = io_decode_csr == 12'hb9e; // @[csr.scala 259:76:Sodor3Stage.fir@2213.4]
  assign _T_637 = io_decode_csr == 12'hb1f; // @[csr.scala 259:76:Sodor3Stage.fir@2214.4]
  assign _T_639 = io_decode_csr == 12'hb9f; // @[csr.scala 259:76:Sodor3Stage.fir@2215.4]
  assign _T_641 = io_decode_csr == 12'hb20; // @[csr.scala 259:76:Sodor3Stage.fir@2216.4]
  assign _T_643 = io_decode_csr == 12'hba0; // @[csr.scala 259:76:Sodor3Stage.fir@2217.4]
  assign _T_645 = io_decode_csr == 12'hb21; // @[csr.scala 259:76:Sodor3Stage.fir@2218.4]
  assign _T_647 = io_decode_csr == 12'hba1; // @[csr.scala 259:76:Sodor3Stage.fir@2219.4]
  assign _T_649 = io_decode_csr == 12'hb22; // @[csr.scala 259:76:Sodor3Stage.fir@2220.4]
  assign _T_651 = io_decode_csr == 12'hba2; // @[csr.scala 259:76:Sodor3Stage.fir@2221.4]
  assign _T_653 = io_decode_csr == 12'hb80; // @[csr.scala 259:76:Sodor3Stage.fir@2222.4]
  assign _T_655 = io_decode_csr == 12'hb82; // @[csr.scala 259:76:Sodor3Stage.fir@2223.4]
  assign _T_656 = io_decode_csr[9:8]; // @[csr.scala 261:57:Sodor3Stage.fir@2224.4]
  assign priv_sufficient = reg_mstatus_prv >= _T_656; // @[csr.scala 261:41:Sodor3Stage.fir@2225.4]
  assign _T_657 = io_decode_csr[11:10]; // @[csr.scala 262:32:Sodor3Stage.fir@2226.4]
  assign _T_658 = ~ _T_657; // @[csr.scala 262:40:Sodor3Stage.fir@2227.4]
  assign read_only = _T_658 == 2'h0; // @[csr.scala 262:40:Sodor3Stage.fir@2228.4]
  assign _T_660 = io_rw_cmd != 3'h5; // @[csr.scala 263:38:Sodor3Stage.fir@2229.4]
  assign _T_661 = cpu_ren & _T_660; // @[csr.scala 263:25:Sodor3Stage.fir@2230.4]
  assign cpu_wen = _T_661 & priv_sufficient; // @[csr.scala 263:47:Sodor3Stage.fir@2231.4]
  assign _T_663 = read_only == 1'h0; // @[csr.scala 264:24:Sodor3Stage.fir@2232.4]
  assign wen = cpu_wen & _T_663; // @[csr.scala 264:21:Sodor3Stage.fir@2233.4]
  assign _T_664 = io_rw_cmd == 3'h2; // @[util.scala 25:47:Sodor3Stage.fir@2234.4]
  assign _T_665 = io_rw_cmd == 3'h3; // @[util.scala 25:47:Sodor3Stage.fir@2235.4]
  assign _T_666 = _T_664 | _T_665; // @[util.scala 25:62:Sodor3Stage.fir@2236.4]
  assign _T_668 = _T_666 ? io_rw_rdata : 32'h0; // @[csr.scala 390:9:Sodor3Stage.fir@2237.4]
  assign _T_669 = _T_668 | io_rw_wdata; // @[csr.scala 390:53:Sodor3Stage.fir@2238.4]
  assign _T_672 = _T_665 ? io_rw_wdata : 32'h0; // @[csr.scala 390:68:Sodor3Stage.fir@2240.4]
  assign _T_673 = ~ _T_672; // @[csr.scala 390:64:Sodor3Stage.fir@2241.4]
  assign wdata = _T_669 & _T_673; // @[csr.scala 390:62:Sodor3Stage.fir@2242.4]
  assign _T_675 = io_decode_csr[2:0]; // @[csr.scala 267:36:Sodor3Stage.fir@2243.4]
  assign opcode = 8'h1 << _T_675; // @[csr.scala 267:20:Sodor3Stage.fir@2244.4]
  assign _T_676 = opcode[0]; // @[csr.scala 268:40:Sodor3Stage.fir@2245.4]
  assign insn_call = system_insn & _T_676; // @[csr.scala 268:31:Sodor3Stage.fir@2246.4]
  assign _T_677 = opcode[1]; // @[csr.scala 269:41:Sodor3Stage.fir@2247.4]
  assign insn_break = system_insn & _T_677; // @[csr.scala 269:32:Sodor3Stage.fir@2248.4]
  assign _T_678 = opcode[2]; // @[csr.scala 270:39:Sodor3Stage.fir@2249.4]
  assign _T_679 = system_insn & _T_678; // @[csr.scala 270:30:Sodor3Stage.fir@2250.4]
  assign insn_ret = _T_679 & priv_sufficient; // @[csr.scala 270:43:Sodor3Stage.fir@2251.4]
  assign _T_962 = insn_call | insn_break; // @[csr.scala 282:24:Sodor3Stage.fir@2469.4]
  assign _GEN_4 = io_exception ? io_pc : reg_mepc; // @[csr.scala 285:23:Sodor3Stage.fir@2472.4]
  assign _T_966 = insn_ret + io_exception; // @[Bitwise.scala 48:55:Sodor3Stage.fir@2477.4]
  assign _T_968 = _T_966 <= 2'h1; // @[csr.scala 291:52:Sodor3Stage.fir@2478.4]
  assign _T_970 = _T_968 | reset; // @[csr.scala 291:9:Sodor3Stage.fir@2480.4]
  assign _T_975 = io_decode_csr[10]; // @[csr.scala 298:33:Sodor3Stage.fir@2490.4]
  assign _T_976 = insn_ret & _T_975; // @[csr.scala 298:17:Sodor3Stage.fir@2491.4]
  assign _GEN_8 = _T_976 ? reg_dpc : 32'h80000004; // @[csr.scala 298:38:Sodor3Stage.fir@2492.4]
  assign _T_980 = _T_975 == 1'h0; // @[csr.scala 305:21:Sodor3Stage.fir@2498.4]
  assign _T_981 = insn_ret & _T_980; // @[csr.scala 305:18:Sodor3Stage.fir@2499.4]
  assign _GEN_12 = _T_981 ? reg_mepc : _GEN_8; // @[csr.scala 305:41:Sodor3Stage.fir@2500.4]
  assign _GEN_390 = {{2'd0}, reg_mstatus_prv}; // @[csr.scala 315:35:Sodor3Stage.fir@2508.6]
  assign _T_985 = _GEN_390 + 4'h8; // @[csr.scala 315:35:Sodor3Stage.fir@2508.6]
  assign _T_986 = _T_985[3:0]; // @[csr.scala 315:35:Sodor3Stage.fir@2509.6]
  assign _GEN_13 = insn_call ? 32'h80000004 : _GEN_12; // @[csr.scala 313:18:Sodor3Stage.fir@2506.4]
  assign _T_991 = _T_487 ? _T_185 : 64'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2518.4]
  assign _T_993 = _T_489 ? _T_197 : 64'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2519.4]
  assign _T_995 = _T_491 ? 16'h8000 : 16'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2520.4]
  assign _T_1001 = _T_497 ? 9'h100 : 9'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2523.4]
  assign _T_1003 = _T_499 ? read_mstatus : 35'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2524.4]
  assign _T_1005 = _T_501 ? 9'h100 : 9'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2525.4]
  assign _T_1007 = _T_503 ? _T_454 : 16'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2526.4]
  assign _T_1009 = _T_505 ? _T_469 : 16'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2527.4]
  assign _T_1011 = _T_507 ? reg_mscratch : 32'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2528.4]
  assign _T_1013 = _T_509 ? reg_mepc : 32'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2529.4]
  assign _T_1015 = _T_511 ? reg_mtval : 32'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2530.4]
  assign _T_1017 = _T_513 ? reg_mcause : 32'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2531.4]
  assign _T_1021 = _T_517 ? _T_483 : 32'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2533.4]
  assign _T_1023 = _T_519 ? reg_dpc : 32'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2534.4]
  assign _T_1025 = _T_521 ? reg_dscratch : 32'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2535.4]
  assign _T_1027 = _T_523 ? reg_medeleg : 32'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2536.4]
  assign _T_1029 = _T_525 ? _T_200 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2537.4]
  assign _T_1031 = _T_527 ? _T_200 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2538.4]
  assign _T_1033 = _T_529 ? _T_203 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2539.4]
  assign _T_1035 = _T_531 ? _T_203 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2540.4]
  assign _T_1037 = _T_533 ? _T_206 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2541.4]
  assign _T_1039 = _T_535 ? _T_206 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2542.4]
  assign _T_1041 = _T_537 ? _T_209 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2543.4]
  assign _T_1043 = _T_539 ? _T_209 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2544.4]
  assign _T_1045 = _T_541 ? _T_212 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2545.4]
  assign _T_1047 = _T_543 ? _T_212 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2546.4]
  assign _T_1049 = _T_545 ? _T_215 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2547.4]
  assign _T_1051 = _T_547 ? _T_215 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2548.4]
  assign _T_1053 = _T_549 ? _T_218 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2549.4]
  assign _T_1055 = _T_551 ? _T_218 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2550.4]
  assign _T_1057 = _T_553 ? _T_221 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2551.4]
  assign _T_1059 = _T_555 ? _T_221 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2552.4]
  assign _T_1061 = _T_557 ? _T_224 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2553.4]
  assign _T_1063 = _T_559 ? _T_224 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2554.4]
  assign _T_1065 = _T_561 ? _T_227 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2555.4]
  assign _T_1067 = _T_563 ? _T_227 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2556.4]
  assign _T_1069 = _T_565 ? _T_230 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2557.4]
  assign _T_1071 = _T_567 ? _T_230 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2558.4]
  assign _T_1073 = _T_569 ? _T_233 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2559.4]
  assign _T_1075 = _T_571 ? _T_233 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2560.4]
  assign _T_1077 = _T_573 ? _T_236 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2561.4]
  assign _T_1079 = _T_575 ? _T_236 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2562.4]
  assign _T_1081 = _T_577 ? _T_239 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2563.4]
  assign _T_1083 = _T_579 ? _T_239 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2564.4]
  assign _T_1085 = _T_581 ? _T_242 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2565.4]
  assign _T_1087 = _T_583 ? _T_242 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2566.4]
  assign _T_1089 = _T_585 ? _T_245 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2567.4]
  assign _T_1091 = _T_587 ? _T_245 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2568.4]
  assign _T_1093 = _T_589 ? _T_248 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2569.4]
  assign _T_1095 = _T_591 ? _T_248 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2570.4]
  assign _T_1097 = _T_593 ? _T_251 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2571.4]
  assign _T_1099 = _T_595 ? _T_251 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2572.4]
  assign _T_1101 = _T_597 ? _T_254 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2573.4]
  assign _T_1103 = _T_599 ? _T_254 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2574.4]
  assign _T_1105 = _T_601 ? _T_257 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2575.4]
  assign _T_1107 = _T_603 ? _T_257 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2576.4]
  assign _T_1109 = _T_605 ? _T_260 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2577.4]
  assign _T_1111 = _T_607 ? _T_260 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2578.4]
  assign _T_1113 = _T_609 ? _T_263 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2579.4]
  assign _T_1115 = _T_611 ? _T_263 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2580.4]
  assign _T_1117 = _T_613 ? _T_266 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2581.4]
  assign _T_1119 = _T_615 ? _T_266 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2582.4]
  assign _T_1121 = _T_617 ? _T_269 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2583.4]
  assign _T_1123 = _T_619 ? _T_269 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2584.4]
  assign _T_1125 = _T_621 ? _T_272 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2585.4]
  assign _T_1127 = _T_623 ? _T_272 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2586.4]
  assign _T_1129 = _T_625 ? _T_275 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2587.4]
  assign _T_1131 = _T_627 ? _T_275 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2588.4]
  assign _T_1133 = _T_629 ? _T_278 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2589.4]
  assign _T_1135 = _T_631 ? _T_278 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2590.4]
  assign _T_1137 = _T_633 ? _T_281 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2591.4]
  assign _T_1139 = _T_635 ? _T_281 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2592.4]
  assign _T_1141 = _T_637 ? _T_284 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2593.4]
  assign _T_1143 = _T_639 ? _T_284 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2594.4]
  assign _T_1145 = _T_641 ? _T_287 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2595.4]
  assign _T_1147 = _T_643 ? _T_287 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2596.4]
  assign _T_1149 = _T_645 ? _T_290 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2597.4]
  assign _T_1151 = _T_647 ? _T_290 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2598.4]
  assign _T_1153 = _T_649 ? _T_293 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2599.4]
  assign _T_1155 = _T_651 ? _T_293 : 40'h0; // @[Mux.scala 19:72:Sodor3Stage.fir@2600.4]
  assign _T_1160 = _T_991 | _T_993; // @[Mux.scala 19:72:Sodor3Stage.fir@2603.4]
  assign _GEN_391 = {{48'd0}, _T_995}; // @[Mux.scala 19:72:Sodor3Stage.fir@2604.4]
  assign _T_1161 = _T_1160 | _GEN_391; // @[Mux.scala 19:72:Sodor3Stage.fir@2604.4]
  assign _GEN_392 = {{55'd0}, _T_1001}; // @[Mux.scala 19:72:Sodor3Stage.fir@2607.4]
  assign _T_1164 = _T_1161 | _GEN_392; // @[Mux.scala 19:72:Sodor3Stage.fir@2607.4]
  assign _GEN_393 = {{29'd0}, _T_1003}; // @[Mux.scala 19:72:Sodor3Stage.fir@2608.4]
  assign _T_1165 = _T_1164 | _GEN_393; // @[Mux.scala 19:72:Sodor3Stage.fir@2608.4]
  assign _GEN_394 = {{55'd0}, _T_1005}; // @[Mux.scala 19:72:Sodor3Stage.fir@2609.4]
  assign _T_1166 = _T_1165 | _GEN_394; // @[Mux.scala 19:72:Sodor3Stage.fir@2609.4]
  assign _GEN_395 = {{48'd0}, _T_1007}; // @[Mux.scala 19:72:Sodor3Stage.fir@2610.4]
  assign _T_1167 = _T_1166 | _GEN_395; // @[Mux.scala 19:72:Sodor3Stage.fir@2610.4]
  assign _GEN_396 = {{48'd0}, _T_1009}; // @[Mux.scala 19:72:Sodor3Stage.fir@2611.4]
  assign _T_1168 = _T_1167 | _GEN_396; // @[Mux.scala 19:72:Sodor3Stage.fir@2611.4]
  assign _GEN_397 = {{32'd0}, _T_1011}; // @[Mux.scala 19:72:Sodor3Stage.fir@2612.4]
  assign _T_1169 = _T_1168 | _GEN_397; // @[Mux.scala 19:72:Sodor3Stage.fir@2612.4]
  assign _GEN_398 = {{32'd0}, _T_1013}; // @[Mux.scala 19:72:Sodor3Stage.fir@2613.4]
  assign _T_1170 = _T_1169 | _GEN_398; // @[Mux.scala 19:72:Sodor3Stage.fir@2613.4]
  assign _GEN_399 = {{32'd0}, _T_1015}; // @[Mux.scala 19:72:Sodor3Stage.fir@2614.4]
  assign _T_1171 = _T_1170 | _GEN_399; // @[Mux.scala 19:72:Sodor3Stage.fir@2614.4]
  assign _GEN_400 = {{32'd0}, _T_1017}; // @[Mux.scala 19:72:Sodor3Stage.fir@2615.4]
  assign _T_1172 = _T_1171 | _GEN_400; // @[Mux.scala 19:72:Sodor3Stage.fir@2615.4]
  assign _GEN_401 = {{32'd0}, _T_1021}; // @[Mux.scala 19:72:Sodor3Stage.fir@2617.4]
  assign _T_1174 = _T_1172 | _GEN_401; // @[Mux.scala 19:72:Sodor3Stage.fir@2617.4]
  assign _GEN_402 = {{32'd0}, _T_1023}; // @[Mux.scala 19:72:Sodor3Stage.fir@2618.4]
  assign _T_1175 = _T_1174 | _GEN_402; // @[Mux.scala 19:72:Sodor3Stage.fir@2618.4]
  assign _GEN_403 = {{32'd0}, _T_1025}; // @[Mux.scala 19:72:Sodor3Stage.fir@2619.4]
  assign _T_1176 = _T_1175 | _GEN_403; // @[Mux.scala 19:72:Sodor3Stage.fir@2619.4]
  assign _GEN_404 = {{32'd0}, _T_1027}; // @[Mux.scala 19:72:Sodor3Stage.fir@2620.4]
  assign _T_1177 = _T_1176 | _GEN_404; // @[Mux.scala 19:72:Sodor3Stage.fir@2620.4]
  assign _GEN_405 = {{24'd0}, _T_1029}; // @[Mux.scala 19:72:Sodor3Stage.fir@2621.4]
  assign _T_1178 = _T_1177 | _GEN_405; // @[Mux.scala 19:72:Sodor3Stage.fir@2621.4]
  assign _GEN_406 = {{24'd0}, _T_1031}; // @[Mux.scala 19:72:Sodor3Stage.fir@2622.4]
  assign _T_1179 = _T_1178 | _GEN_406; // @[Mux.scala 19:72:Sodor3Stage.fir@2622.4]
  assign _GEN_407 = {{24'd0}, _T_1033}; // @[Mux.scala 19:72:Sodor3Stage.fir@2623.4]
  assign _T_1180 = _T_1179 | _GEN_407; // @[Mux.scala 19:72:Sodor3Stage.fir@2623.4]
  assign _GEN_408 = {{24'd0}, _T_1035}; // @[Mux.scala 19:72:Sodor3Stage.fir@2624.4]
  assign _T_1181 = _T_1180 | _GEN_408; // @[Mux.scala 19:72:Sodor3Stage.fir@2624.4]
  assign _GEN_409 = {{24'd0}, _T_1037}; // @[Mux.scala 19:72:Sodor3Stage.fir@2625.4]
  assign _T_1182 = _T_1181 | _GEN_409; // @[Mux.scala 19:72:Sodor3Stage.fir@2625.4]
  assign _GEN_410 = {{24'd0}, _T_1039}; // @[Mux.scala 19:72:Sodor3Stage.fir@2626.4]
  assign _T_1183 = _T_1182 | _GEN_410; // @[Mux.scala 19:72:Sodor3Stage.fir@2626.4]
  assign _GEN_411 = {{24'd0}, _T_1041}; // @[Mux.scala 19:72:Sodor3Stage.fir@2627.4]
  assign _T_1184 = _T_1183 | _GEN_411; // @[Mux.scala 19:72:Sodor3Stage.fir@2627.4]
  assign _GEN_412 = {{24'd0}, _T_1043}; // @[Mux.scala 19:72:Sodor3Stage.fir@2628.4]
  assign _T_1185 = _T_1184 | _GEN_412; // @[Mux.scala 19:72:Sodor3Stage.fir@2628.4]
  assign _GEN_413 = {{24'd0}, _T_1045}; // @[Mux.scala 19:72:Sodor3Stage.fir@2629.4]
  assign _T_1186 = _T_1185 | _GEN_413; // @[Mux.scala 19:72:Sodor3Stage.fir@2629.4]
  assign _GEN_414 = {{24'd0}, _T_1047}; // @[Mux.scala 19:72:Sodor3Stage.fir@2630.4]
  assign _T_1187 = _T_1186 | _GEN_414; // @[Mux.scala 19:72:Sodor3Stage.fir@2630.4]
  assign _GEN_415 = {{24'd0}, _T_1049}; // @[Mux.scala 19:72:Sodor3Stage.fir@2631.4]
  assign _T_1188 = _T_1187 | _GEN_415; // @[Mux.scala 19:72:Sodor3Stage.fir@2631.4]
  assign _GEN_416 = {{24'd0}, _T_1051}; // @[Mux.scala 19:72:Sodor3Stage.fir@2632.4]
  assign _T_1189 = _T_1188 | _GEN_416; // @[Mux.scala 19:72:Sodor3Stage.fir@2632.4]
  assign _GEN_417 = {{24'd0}, _T_1053}; // @[Mux.scala 19:72:Sodor3Stage.fir@2633.4]
  assign _T_1190 = _T_1189 | _GEN_417; // @[Mux.scala 19:72:Sodor3Stage.fir@2633.4]
  assign _GEN_418 = {{24'd0}, _T_1055}; // @[Mux.scala 19:72:Sodor3Stage.fir@2634.4]
  assign _T_1191 = _T_1190 | _GEN_418; // @[Mux.scala 19:72:Sodor3Stage.fir@2634.4]
  assign _GEN_419 = {{24'd0}, _T_1057}; // @[Mux.scala 19:72:Sodor3Stage.fir@2635.4]
  assign _T_1192 = _T_1191 | _GEN_419; // @[Mux.scala 19:72:Sodor3Stage.fir@2635.4]
  assign _GEN_420 = {{24'd0}, _T_1059}; // @[Mux.scala 19:72:Sodor3Stage.fir@2636.4]
  assign _T_1193 = _T_1192 | _GEN_420; // @[Mux.scala 19:72:Sodor3Stage.fir@2636.4]
  assign _GEN_421 = {{24'd0}, _T_1061}; // @[Mux.scala 19:72:Sodor3Stage.fir@2637.4]
  assign _T_1194 = _T_1193 | _GEN_421; // @[Mux.scala 19:72:Sodor3Stage.fir@2637.4]
  assign _GEN_422 = {{24'd0}, _T_1063}; // @[Mux.scala 19:72:Sodor3Stage.fir@2638.4]
  assign _T_1195 = _T_1194 | _GEN_422; // @[Mux.scala 19:72:Sodor3Stage.fir@2638.4]
  assign _GEN_423 = {{24'd0}, _T_1065}; // @[Mux.scala 19:72:Sodor3Stage.fir@2639.4]
  assign _T_1196 = _T_1195 | _GEN_423; // @[Mux.scala 19:72:Sodor3Stage.fir@2639.4]
  assign _GEN_424 = {{24'd0}, _T_1067}; // @[Mux.scala 19:72:Sodor3Stage.fir@2640.4]
  assign _T_1197 = _T_1196 | _GEN_424; // @[Mux.scala 19:72:Sodor3Stage.fir@2640.4]
  assign _GEN_425 = {{24'd0}, _T_1069}; // @[Mux.scala 19:72:Sodor3Stage.fir@2641.4]
  assign _T_1198 = _T_1197 | _GEN_425; // @[Mux.scala 19:72:Sodor3Stage.fir@2641.4]
  assign _GEN_426 = {{24'd0}, _T_1071}; // @[Mux.scala 19:72:Sodor3Stage.fir@2642.4]
  assign _T_1199 = _T_1198 | _GEN_426; // @[Mux.scala 19:72:Sodor3Stage.fir@2642.4]
  assign _GEN_427 = {{24'd0}, _T_1073}; // @[Mux.scala 19:72:Sodor3Stage.fir@2643.4]
  assign _T_1200 = _T_1199 | _GEN_427; // @[Mux.scala 19:72:Sodor3Stage.fir@2643.4]
  assign _GEN_428 = {{24'd0}, _T_1075}; // @[Mux.scala 19:72:Sodor3Stage.fir@2644.4]
  assign _T_1201 = _T_1200 | _GEN_428; // @[Mux.scala 19:72:Sodor3Stage.fir@2644.4]
  assign _GEN_429 = {{24'd0}, _T_1077}; // @[Mux.scala 19:72:Sodor3Stage.fir@2645.4]
  assign _T_1202 = _T_1201 | _GEN_429; // @[Mux.scala 19:72:Sodor3Stage.fir@2645.4]
  assign _GEN_430 = {{24'd0}, _T_1079}; // @[Mux.scala 19:72:Sodor3Stage.fir@2646.4]
  assign _T_1203 = _T_1202 | _GEN_430; // @[Mux.scala 19:72:Sodor3Stage.fir@2646.4]
  assign _GEN_431 = {{24'd0}, _T_1081}; // @[Mux.scala 19:72:Sodor3Stage.fir@2647.4]
  assign _T_1204 = _T_1203 | _GEN_431; // @[Mux.scala 19:72:Sodor3Stage.fir@2647.4]
  assign _GEN_432 = {{24'd0}, _T_1083}; // @[Mux.scala 19:72:Sodor3Stage.fir@2648.4]
  assign _T_1205 = _T_1204 | _GEN_432; // @[Mux.scala 19:72:Sodor3Stage.fir@2648.4]
  assign _GEN_433 = {{24'd0}, _T_1085}; // @[Mux.scala 19:72:Sodor3Stage.fir@2649.4]
  assign _T_1206 = _T_1205 | _GEN_433; // @[Mux.scala 19:72:Sodor3Stage.fir@2649.4]
  assign _GEN_434 = {{24'd0}, _T_1087}; // @[Mux.scala 19:72:Sodor3Stage.fir@2650.4]
  assign _T_1207 = _T_1206 | _GEN_434; // @[Mux.scala 19:72:Sodor3Stage.fir@2650.4]
  assign _GEN_435 = {{24'd0}, _T_1089}; // @[Mux.scala 19:72:Sodor3Stage.fir@2651.4]
  assign _T_1208 = _T_1207 | _GEN_435; // @[Mux.scala 19:72:Sodor3Stage.fir@2651.4]
  assign _GEN_436 = {{24'd0}, _T_1091}; // @[Mux.scala 19:72:Sodor3Stage.fir@2652.4]
  assign _T_1209 = _T_1208 | _GEN_436; // @[Mux.scala 19:72:Sodor3Stage.fir@2652.4]
  assign _GEN_437 = {{24'd0}, _T_1093}; // @[Mux.scala 19:72:Sodor3Stage.fir@2653.4]
  assign _T_1210 = _T_1209 | _GEN_437; // @[Mux.scala 19:72:Sodor3Stage.fir@2653.4]
  assign _GEN_438 = {{24'd0}, _T_1095}; // @[Mux.scala 19:72:Sodor3Stage.fir@2654.4]
  assign _T_1211 = _T_1210 | _GEN_438; // @[Mux.scala 19:72:Sodor3Stage.fir@2654.4]
  assign _GEN_439 = {{24'd0}, _T_1097}; // @[Mux.scala 19:72:Sodor3Stage.fir@2655.4]
  assign _T_1212 = _T_1211 | _GEN_439; // @[Mux.scala 19:72:Sodor3Stage.fir@2655.4]
  assign _GEN_440 = {{24'd0}, _T_1099}; // @[Mux.scala 19:72:Sodor3Stage.fir@2656.4]
  assign _T_1213 = _T_1212 | _GEN_440; // @[Mux.scala 19:72:Sodor3Stage.fir@2656.4]
  assign _GEN_441 = {{24'd0}, _T_1101}; // @[Mux.scala 19:72:Sodor3Stage.fir@2657.4]
  assign _T_1214 = _T_1213 | _GEN_441; // @[Mux.scala 19:72:Sodor3Stage.fir@2657.4]
  assign _GEN_442 = {{24'd0}, _T_1103}; // @[Mux.scala 19:72:Sodor3Stage.fir@2658.4]
  assign _T_1215 = _T_1214 | _GEN_442; // @[Mux.scala 19:72:Sodor3Stage.fir@2658.4]
  assign _GEN_443 = {{24'd0}, _T_1105}; // @[Mux.scala 19:72:Sodor3Stage.fir@2659.4]
  assign _T_1216 = _T_1215 | _GEN_443; // @[Mux.scala 19:72:Sodor3Stage.fir@2659.4]
  assign _GEN_444 = {{24'd0}, _T_1107}; // @[Mux.scala 19:72:Sodor3Stage.fir@2660.4]
  assign _T_1217 = _T_1216 | _GEN_444; // @[Mux.scala 19:72:Sodor3Stage.fir@2660.4]
  assign _GEN_445 = {{24'd0}, _T_1109}; // @[Mux.scala 19:72:Sodor3Stage.fir@2661.4]
  assign _T_1218 = _T_1217 | _GEN_445; // @[Mux.scala 19:72:Sodor3Stage.fir@2661.4]
  assign _GEN_446 = {{24'd0}, _T_1111}; // @[Mux.scala 19:72:Sodor3Stage.fir@2662.4]
  assign _T_1219 = _T_1218 | _GEN_446; // @[Mux.scala 19:72:Sodor3Stage.fir@2662.4]
  assign _GEN_447 = {{24'd0}, _T_1113}; // @[Mux.scala 19:72:Sodor3Stage.fir@2663.4]
  assign _T_1220 = _T_1219 | _GEN_447; // @[Mux.scala 19:72:Sodor3Stage.fir@2663.4]
  assign _GEN_448 = {{24'd0}, _T_1115}; // @[Mux.scala 19:72:Sodor3Stage.fir@2664.4]
  assign _T_1221 = _T_1220 | _GEN_448; // @[Mux.scala 19:72:Sodor3Stage.fir@2664.4]
  assign _GEN_449 = {{24'd0}, _T_1117}; // @[Mux.scala 19:72:Sodor3Stage.fir@2665.4]
  assign _T_1222 = _T_1221 | _GEN_449; // @[Mux.scala 19:72:Sodor3Stage.fir@2665.4]
  assign _GEN_450 = {{24'd0}, _T_1119}; // @[Mux.scala 19:72:Sodor3Stage.fir@2666.4]
  assign _T_1223 = _T_1222 | _GEN_450; // @[Mux.scala 19:72:Sodor3Stage.fir@2666.4]
  assign _GEN_451 = {{24'd0}, _T_1121}; // @[Mux.scala 19:72:Sodor3Stage.fir@2667.4]
  assign _T_1224 = _T_1223 | _GEN_451; // @[Mux.scala 19:72:Sodor3Stage.fir@2667.4]
  assign _GEN_452 = {{24'd0}, _T_1123}; // @[Mux.scala 19:72:Sodor3Stage.fir@2668.4]
  assign _T_1225 = _T_1224 | _GEN_452; // @[Mux.scala 19:72:Sodor3Stage.fir@2668.4]
  assign _GEN_453 = {{24'd0}, _T_1125}; // @[Mux.scala 19:72:Sodor3Stage.fir@2669.4]
  assign _T_1226 = _T_1225 | _GEN_453; // @[Mux.scala 19:72:Sodor3Stage.fir@2669.4]
  assign _GEN_454 = {{24'd0}, _T_1127}; // @[Mux.scala 19:72:Sodor3Stage.fir@2670.4]
  assign _T_1227 = _T_1226 | _GEN_454; // @[Mux.scala 19:72:Sodor3Stage.fir@2670.4]
  assign _GEN_455 = {{24'd0}, _T_1129}; // @[Mux.scala 19:72:Sodor3Stage.fir@2671.4]
  assign _T_1228 = _T_1227 | _GEN_455; // @[Mux.scala 19:72:Sodor3Stage.fir@2671.4]
  assign _GEN_456 = {{24'd0}, _T_1131}; // @[Mux.scala 19:72:Sodor3Stage.fir@2672.4]
  assign _T_1229 = _T_1228 | _GEN_456; // @[Mux.scala 19:72:Sodor3Stage.fir@2672.4]
  assign _GEN_457 = {{24'd0}, _T_1133}; // @[Mux.scala 19:72:Sodor3Stage.fir@2673.4]
  assign _T_1230 = _T_1229 | _GEN_457; // @[Mux.scala 19:72:Sodor3Stage.fir@2673.4]
  assign _GEN_458 = {{24'd0}, _T_1135}; // @[Mux.scala 19:72:Sodor3Stage.fir@2674.4]
  assign _T_1231 = _T_1230 | _GEN_458; // @[Mux.scala 19:72:Sodor3Stage.fir@2674.4]
  assign _GEN_459 = {{24'd0}, _T_1137}; // @[Mux.scala 19:72:Sodor3Stage.fir@2675.4]
  assign _T_1232 = _T_1231 | _GEN_459; // @[Mux.scala 19:72:Sodor3Stage.fir@2675.4]
  assign _GEN_460 = {{24'd0}, _T_1139}; // @[Mux.scala 19:72:Sodor3Stage.fir@2676.4]
  assign _T_1233 = _T_1232 | _GEN_460; // @[Mux.scala 19:72:Sodor3Stage.fir@2676.4]
  assign _GEN_461 = {{24'd0}, _T_1141}; // @[Mux.scala 19:72:Sodor3Stage.fir@2677.4]
  assign _T_1234 = _T_1233 | _GEN_461; // @[Mux.scala 19:72:Sodor3Stage.fir@2677.4]
  assign _GEN_462 = {{24'd0}, _T_1143}; // @[Mux.scala 19:72:Sodor3Stage.fir@2678.4]
  assign _T_1235 = _T_1234 | _GEN_462; // @[Mux.scala 19:72:Sodor3Stage.fir@2678.4]
  assign _GEN_463 = {{24'd0}, _T_1145}; // @[Mux.scala 19:72:Sodor3Stage.fir@2679.4]
  assign _T_1236 = _T_1235 | _GEN_463; // @[Mux.scala 19:72:Sodor3Stage.fir@2679.4]
  assign _GEN_464 = {{24'd0}, _T_1147}; // @[Mux.scala 19:72:Sodor3Stage.fir@2680.4]
  assign _T_1237 = _T_1236 | _GEN_464; // @[Mux.scala 19:72:Sodor3Stage.fir@2680.4]
  assign _GEN_465 = {{24'd0}, _T_1149}; // @[Mux.scala 19:72:Sodor3Stage.fir@2681.4]
  assign _T_1238 = _T_1237 | _GEN_465; // @[Mux.scala 19:72:Sodor3Stage.fir@2681.4]
  assign _GEN_466 = {{24'd0}, _T_1151}; // @[Mux.scala 19:72:Sodor3Stage.fir@2682.4]
  assign _T_1239 = _T_1238 | _GEN_466; // @[Mux.scala 19:72:Sodor3Stage.fir@2682.4]
  assign _GEN_467 = {{24'd0}, _T_1153}; // @[Mux.scala 19:72:Sodor3Stage.fir@2683.4]
  assign _T_1240 = _T_1239 | _GEN_467; // @[Mux.scala 19:72:Sodor3Stage.fir@2683.4]
  assign _GEN_468 = {{24'd0}, _T_1155}; // @[Mux.scala 19:72:Sodor3Stage.fir@2684.4]
  assign _T_1241 = _T_1240 | _GEN_468; // @[Mux.scala 19:72:Sodor3Stage.fir@2684.4]
  assign _T_1252 = wdata[2]; // @[csr.scala 334:43:Sodor3Stage.fir@2697.8]
  assign _T_1262 = wdata[15]; // @[csr.scala 334:43:Sodor3Stage.fir@2717.8]
  assign _T_1270 = {{3'd0}, wdata}; // @[:Sodor3Stage.fir@2730.8]
  assign _T_1274 = _T_1270[3]; // @[csr.scala 341:47:Sodor3Stage.fir@2738.8]
  assign _T_1278 = _T_1270[7]; // @[csr.scala 341:47:Sodor3Stage.fir@2746.8]
  assign _T_1298 = wdata[15:0]; // @[:Sodor3Stage.fir@2783.8]
  assign _T_1302 = _T_1298[3]; // @[csr.scala 346:39:Sodor3Stage.fir@2791.8]
  assign _T_1306 = _T_1298[7]; // @[csr.scala 346:39:Sodor3Stage.fir@2799.8]
  assign _T_1336 = wdata[7:0]; // @[csr.scala 386:47:Sodor3Stage.fir@2859.8]
  assign _T_1337 = _T_200[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@2860.8]
  assign _T_1338 = {_T_1336,_T_1337}; // @[Cat.scala 30:58:Sodor3Stage.fir@2861.8]
  assign _GEN_24 = _T_527 ? {{1'd0}, _T_1338} : _T_201; // @[csr.scala 386:29:Sodor3Stage.fir@2858.6]
  assign _T_1339 = _T_200[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@2865.8]
  assign _T_1340 = {_T_1339,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@2866.8]
  assign _GEN_25 = _T_525 ? {{1'd0}, _T_1340} : _GEN_24; // @[csr.scala 387:29:Sodor3Stage.fir@2864.6]
  assign _T_1342 = _T_203[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@2871.8]
  assign _T_1343 = {_T_1336,_T_1342}; // @[Cat.scala 30:58:Sodor3Stage.fir@2872.8]
  assign _GEN_26 = _T_531 ? {{1'd0}, _T_1343} : _T_204; // @[csr.scala 386:29:Sodor3Stage.fir@2869.6]
  assign _T_1344 = _T_203[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@2876.8]
  assign _T_1345 = {_T_1344,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@2877.8]
  assign _GEN_27 = _T_529 ? {{1'd0}, _T_1345} : _GEN_26; // @[csr.scala 387:29:Sodor3Stage.fir@2875.6]
  assign _T_1347 = _T_206[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@2882.8]
  assign _T_1348 = {_T_1336,_T_1347}; // @[Cat.scala 30:58:Sodor3Stage.fir@2883.8]
  assign _GEN_28 = _T_535 ? {{1'd0}, _T_1348} : _T_207; // @[csr.scala 386:29:Sodor3Stage.fir@2880.6]
  assign _T_1349 = _T_206[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@2887.8]
  assign _T_1350 = {_T_1349,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@2888.8]
  assign _GEN_29 = _T_533 ? {{1'd0}, _T_1350} : _GEN_28; // @[csr.scala 387:29:Sodor3Stage.fir@2886.6]
  assign _T_1352 = _T_209[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@2893.8]
  assign _T_1353 = {_T_1336,_T_1352}; // @[Cat.scala 30:58:Sodor3Stage.fir@2894.8]
  assign _GEN_30 = _T_539 ? {{1'd0}, _T_1353} : _T_210; // @[csr.scala 386:29:Sodor3Stage.fir@2891.6]
  assign _T_1354 = _T_209[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@2898.8]
  assign _T_1355 = {_T_1354,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@2899.8]
  assign _GEN_31 = _T_537 ? {{1'd0}, _T_1355} : _GEN_30; // @[csr.scala 387:29:Sodor3Stage.fir@2897.6]
  assign _T_1357 = _T_212[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@2904.8]
  assign _T_1358 = {_T_1336,_T_1357}; // @[Cat.scala 30:58:Sodor3Stage.fir@2905.8]
  assign _GEN_32 = _T_543 ? {{1'd0}, _T_1358} : _T_213; // @[csr.scala 386:29:Sodor3Stage.fir@2902.6]
  assign _T_1359 = _T_212[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@2909.8]
  assign _T_1360 = {_T_1359,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@2910.8]
  assign _GEN_33 = _T_541 ? {{1'd0}, _T_1360} : _GEN_32; // @[csr.scala 387:29:Sodor3Stage.fir@2908.6]
  assign _T_1362 = _T_215[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@2915.8]
  assign _T_1363 = {_T_1336,_T_1362}; // @[Cat.scala 30:58:Sodor3Stage.fir@2916.8]
  assign _GEN_34 = _T_547 ? {{1'd0}, _T_1363} : _T_216; // @[csr.scala 386:29:Sodor3Stage.fir@2913.6]
  assign _T_1364 = _T_215[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@2920.8]
  assign _T_1365 = {_T_1364,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@2921.8]
  assign _GEN_35 = _T_545 ? {{1'd0}, _T_1365} : _GEN_34; // @[csr.scala 387:29:Sodor3Stage.fir@2919.6]
  assign _T_1367 = _T_218[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@2926.8]
  assign _T_1368 = {_T_1336,_T_1367}; // @[Cat.scala 30:58:Sodor3Stage.fir@2927.8]
  assign _GEN_36 = _T_551 ? {{1'd0}, _T_1368} : _T_219; // @[csr.scala 386:29:Sodor3Stage.fir@2924.6]
  assign _T_1369 = _T_218[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@2931.8]
  assign _T_1370 = {_T_1369,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@2932.8]
  assign _GEN_37 = _T_549 ? {{1'd0}, _T_1370} : _GEN_36; // @[csr.scala 387:29:Sodor3Stage.fir@2930.6]
  assign _T_1372 = _T_221[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@2937.8]
  assign _T_1373 = {_T_1336,_T_1372}; // @[Cat.scala 30:58:Sodor3Stage.fir@2938.8]
  assign _GEN_38 = _T_555 ? {{1'd0}, _T_1373} : _T_222; // @[csr.scala 386:29:Sodor3Stage.fir@2935.6]
  assign _T_1374 = _T_221[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@2942.8]
  assign _T_1375 = {_T_1374,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@2943.8]
  assign _GEN_39 = _T_553 ? {{1'd0}, _T_1375} : _GEN_38; // @[csr.scala 387:29:Sodor3Stage.fir@2941.6]
  assign _T_1377 = _T_224[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@2948.8]
  assign _T_1378 = {_T_1336,_T_1377}; // @[Cat.scala 30:58:Sodor3Stage.fir@2949.8]
  assign _GEN_40 = _T_559 ? {{1'd0}, _T_1378} : _T_225; // @[csr.scala 386:29:Sodor3Stage.fir@2946.6]
  assign _T_1379 = _T_224[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@2953.8]
  assign _T_1380 = {_T_1379,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@2954.8]
  assign _GEN_41 = _T_557 ? {{1'd0}, _T_1380} : _GEN_40; // @[csr.scala 387:29:Sodor3Stage.fir@2952.6]
  assign _T_1382 = _T_227[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@2959.8]
  assign _T_1383 = {_T_1336,_T_1382}; // @[Cat.scala 30:58:Sodor3Stage.fir@2960.8]
  assign _GEN_42 = _T_563 ? {{1'd0}, _T_1383} : _T_228; // @[csr.scala 386:29:Sodor3Stage.fir@2957.6]
  assign _T_1384 = _T_227[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@2964.8]
  assign _T_1385 = {_T_1384,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@2965.8]
  assign _GEN_43 = _T_561 ? {{1'd0}, _T_1385} : _GEN_42; // @[csr.scala 387:29:Sodor3Stage.fir@2963.6]
  assign _T_1387 = _T_230[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@2970.8]
  assign _T_1388 = {_T_1336,_T_1387}; // @[Cat.scala 30:58:Sodor3Stage.fir@2971.8]
  assign _GEN_44 = _T_567 ? {{1'd0}, _T_1388} : _T_231; // @[csr.scala 386:29:Sodor3Stage.fir@2968.6]
  assign _T_1389 = _T_230[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@2975.8]
  assign _T_1390 = {_T_1389,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@2976.8]
  assign _GEN_45 = _T_565 ? {{1'd0}, _T_1390} : _GEN_44; // @[csr.scala 387:29:Sodor3Stage.fir@2974.6]
  assign _T_1392 = _T_233[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@2981.8]
  assign _T_1393 = {_T_1336,_T_1392}; // @[Cat.scala 30:58:Sodor3Stage.fir@2982.8]
  assign _GEN_46 = _T_571 ? {{1'd0}, _T_1393} : _T_234; // @[csr.scala 386:29:Sodor3Stage.fir@2979.6]
  assign _T_1394 = _T_233[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@2986.8]
  assign _T_1395 = {_T_1394,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@2987.8]
  assign _GEN_47 = _T_569 ? {{1'd0}, _T_1395} : _GEN_46; // @[csr.scala 387:29:Sodor3Stage.fir@2985.6]
  assign _T_1397 = _T_236[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@2992.8]
  assign _T_1398 = {_T_1336,_T_1397}; // @[Cat.scala 30:58:Sodor3Stage.fir@2993.8]
  assign _GEN_48 = _T_575 ? {{1'd0}, _T_1398} : _T_237; // @[csr.scala 386:29:Sodor3Stage.fir@2990.6]
  assign _T_1399 = _T_236[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@2997.8]
  assign _T_1400 = {_T_1399,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@2998.8]
  assign _GEN_49 = _T_573 ? {{1'd0}, _T_1400} : _GEN_48; // @[csr.scala 387:29:Sodor3Stage.fir@2996.6]
  assign _T_1402 = _T_239[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@3003.8]
  assign _T_1403 = {_T_1336,_T_1402}; // @[Cat.scala 30:58:Sodor3Stage.fir@3004.8]
  assign _GEN_50 = _T_579 ? {{1'd0}, _T_1403} : _T_240; // @[csr.scala 386:29:Sodor3Stage.fir@3001.6]
  assign _T_1404 = _T_239[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@3008.8]
  assign _T_1405 = {_T_1404,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@3009.8]
  assign _GEN_51 = _T_577 ? {{1'd0}, _T_1405} : _GEN_50; // @[csr.scala 387:29:Sodor3Stage.fir@3007.6]
  assign _T_1407 = _T_242[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@3014.8]
  assign _T_1408 = {_T_1336,_T_1407}; // @[Cat.scala 30:58:Sodor3Stage.fir@3015.8]
  assign _GEN_52 = _T_583 ? {{1'd0}, _T_1408} : _T_243; // @[csr.scala 386:29:Sodor3Stage.fir@3012.6]
  assign _T_1409 = _T_242[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@3019.8]
  assign _T_1410 = {_T_1409,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@3020.8]
  assign _GEN_53 = _T_581 ? {{1'd0}, _T_1410} : _GEN_52; // @[csr.scala 387:29:Sodor3Stage.fir@3018.6]
  assign _T_1412 = _T_245[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@3025.8]
  assign _T_1413 = {_T_1336,_T_1412}; // @[Cat.scala 30:58:Sodor3Stage.fir@3026.8]
  assign _GEN_54 = _T_587 ? {{1'd0}, _T_1413} : _T_246; // @[csr.scala 386:29:Sodor3Stage.fir@3023.6]
  assign _T_1414 = _T_245[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@3030.8]
  assign _T_1415 = {_T_1414,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@3031.8]
  assign _GEN_55 = _T_585 ? {{1'd0}, _T_1415} : _GEN_54; // @[csr.scala 387:29:Sodor3Stage.fir@3029.6]
  assign _T_1417 = _T_248[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@3036.8]
  assign _T_1418 = {_T_1336,_T_1417}; // @[Cat.scala 30:58:Sodor3Stage.fir@3037.8]
  assign _GEN_56 = _T_591 ? {{1'd0}, _T_1418} : _T_249; // @[csr.scala 386:29:Sodor3Stage.fir@3034.6]
  assign _T_1419 = _T_248[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@3041.8]
  assign _T_1420 = {_T_1419,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@3042.8]
  assign _GEN_57 = _T_589 ? {{1'd0}, _T_1420} : _GEN_56; // @[csr.scala 387:29:Sodor3Stage.fir@3040.6]
  assign _T_1422 = _T_251[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@3047.8]
  assign _T_1423 = {_T_1336,_T_1422}; // @[Cat.scala 30:58:Sodor3Stage.fir@3048.8]
  assign _GEN_58 = _T_595 ? {{1'd0}, _T_1423} : _T_252; // @[csr.scala 386:29:Sodor3Stage.fir@3045.6]
  assign _T_1424 = _T_251[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@3052.8]
  assign _T_1425 = {_T_1424,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@3053.8]
  assign _GEN_59 = _T_593 ? {{1'd0}, _T_1425} : _GEN_58; // @[csr.scala 387:29:Sodor3Stage.fir@3051.6]
  assign _T_1427 = _T_254[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@3058.8]
  assign _T_1428 = {_T_1336,_T_1427}; // @[Cat.scala 30:58:Sodor3Stage.fir@3059.8]
  assign _GEN_60 = _T_599 ? {{1'd0}, _T_1428} : _T_255; // @[csr.scala 386:29:Sodor3Stage.fir@3056.6]
  assign _T_1429 = _T_254[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@3063.8]
  assign _T_1430 = {_T_1429,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@3064.8]
  assign _GEN_61 = _T_597 ? {{1'd0}, _T_1430} : _GEN_60; // @[csr.scala 387:29:Sodor3Stage.fir@3062.6]
  assign _T_1432 = _T_257[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@3069.8]
  assign _T_1433 = {_T_1336,_T_1432}; // @[Cat.scala 30:58:Sodor3Stage.fir@3070.8]
  assign _GEN_62 = _T_603 ? {{1'd0}, _T_1433} : _T_258; // @[csr.scala 386:29:Sodor3Stage.fir@3067.6]
  assign _T_1434 = _T_257[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@3074.8]
  assign _T_1435 = {_T_1434,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@3075.8]
  assign _GEN_63 = _T_601 ? {{1'd0}, _T_1435} : _GEN_62; // @[csr.scala 387:29:Sodor3Stage.fir@3073.6]
  assign _T_1437 = _T_260[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@3080.8]
  assign _T_1438 = {_T_1336,_T_1437}; // @[Cat.scala 30:58:Sodor3Stage.fir@3081.8]
  assign _GEN_64 = _T_607 ? {{1'd0}, _T_1438} : _T_261; // @[csr.scala 386:29:Sodor3Stage.fir@3078.6]
  assign _T_1439 = _T_260[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@3085.8]
  assign _T_1440 = {_T_1439,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@3086.8]
  assign _GEN_65 = _T_605 ? {{1'd0}, _T_1440} : _GEN_64; // @[csr.scala 387:29:Sodor3Stage.fir@3084.6]
  assign _T_1442 = _T_263[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@3091.8]
  assign _T_1443 = {_T_1336,_T_1442}; // @[Cat.scala 30:58:Sodor3Stage.fir@3092.8]
  assign _GEN_66 = _T_611 ? {{1'd0}, _T_1443} : _T_264; // @[csr.scala 386:29:Sodor3Stage.fir@3089.6]
  assign _T_1444 = _T_263[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@3096.8]
  assign _T_1445 = {_T_1444,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@3097.8]
  assign _GEN_67 = _T_609 ? {{1'd0}, _T_1445} : _GEN_66; // @[csr.scala 387:29:Sodor3Stage.fir@3095.6]
  assign _T_1447 = _T_266[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@3102.8]
  assign _T_1448 = {_T_1336,_T_1447}; // @[Cat.scala 30:58:Sodor3Stage.fir@3103.8]
  assign _GEN_68 = _T_615 ? {{1'd0}, _T_1448} : _T_267; // @[csr.scala 386:29:Sodor3Stage.fir@3100.6]
  assign _T_1449 = _T_266[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@3107.8]
  assign _T_1450 = {_T_1449,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@3108.8]
  assign _GEN_69 = _T_613 ? {{1'd0}, _T_1450} : _GEN_68; // @[csr.scala 387:29:Sodor3Stage.fir@3106.6]
  assign _T_1452 = _T_269[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@3113.8]
  assign _T_1453 = {_T_1336,_T_1452}; // @[Cat.scala 30:58:Sodor3Stage.fir@3114.8]
  assign _GEN_70 = _T_619 ? {{1'd0}, _T_1453} : _T_270; // @[csr.scala 386:29:Sodor3Stage.fir@3111.6]
  assign _T_1454 = _T_269[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@3118.8]
  assign _T_1455 = {_T_1454,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@3119.8]
  assign _GEN_71 = _T_617 ? {{1'd0}, _T_1455} : _GEN_70; // @[csr.scala 387:29:Sodor3Stage.fir@3117.6]
  assign _T_1457 = _T_272[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@3124.8]
  assign _T_1458 = {_T_1336,_T_1457}; // @[Cat.scala 30:58:Sodor3Stage.fir@3125.8]
  assign _GEN_72 = _T_623 ? {{1'd0}, _T_1458} : _T_273; // @[csr.scala 386:29:Sodor3Stage.fir@3122.6]
  assign _T_1459 = _T_272[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@3129.8]
  assign _T_1460 = {_T_1459,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@3130.8]
  assign _GEN_73 = _T_621 ? {{1'd0}, _T_1460} : _GEN_72; // @[csr.scala 387:29:Sodor3Stage.fir@3128.6]
  assign _T_1462 = _T_275[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@3135.8]
  assign _T_1463 = {_T_1336,_T_1462}; // @[Cat.scala 30:58:Sodor3Stage.fir@3136.8]
  assign _GEN_74 = _T_627 ? {{1'd0}, _T_1463} : _T_276; // @[csr.scala 386:29:Sodor3Stage.fir@3133.6]
  assign _T_1464 = _T_275[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@3140.8]
  assign _T_1465 = {_T_1464,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@3141.8]
  assign _GEN_75 = _T_625 ? {{1'd0}, _T_1465} : _GEN_74; // @[csr.scala 387:29:Sodor3Stage.fir@3139.6]
  assign _T_1467 = _T_278[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@3146.8]
  assign _T_1468 = {_T_1336,_T_1467}; // @[Cat.scala 30:58:Sodor3Stage.fir@3147.8]
  assign _GEN_76 = _T_631 ? {{1'd0}, _T_1468} : _T_279; // @[csr.scala 386:29:Sodor3Stage.fir@3144.6]
  assign _T_1469 = _T_278[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@3151.8]
  assign _T_1470 = {_T_1469,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@3152.8]
  assign _GEN_77 = _T_629 ? {{1'd0}, _T_1470} : _GEN_76; // @[csr.scala 387:29:Sodor3Stage.fir@3150.6]
  assign _T_1472 = _T_281[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@3157.8]
  assign _T_1473 = {_T_1336,_T_1472}; // @[Cat.scala 30:58:Sodor3Stage.fir@3158.8]
  assign _GEN_78 = _T_635 ? {{1'd0}, _T_1473} : _T_282; // @[csr.scala 386:29:Sodor3Stage.fir@3155.6]
  assign _T_1474 = _T_281[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@3162.8]
  assign _T_1475 = {_T_1474,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@3163.8]
  assign _GEN_79 = _T_633 ? {{1'd0}, _T_1475} : _GEN_78; // @[csr.scala 387:29:Sodor3Stage.fir@3161.6]
  assign _T_1477 = _T_284[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@3168.8]
  assign _T_1478 = {_T_1336,_T_1477}; // @[Cat.scala 30:58:Sodor3Stage.fir@3169.8]
  assign _GEN_80 = _T_639 ? {{1'd0}, _T_1478} : _T_285; // @[csr.scala 386:29:Sodor3Stage.fir@3166.6]
  assign _T_1479 = _T_284[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@3173.8]
  assign _T_1480 = {_T_1479,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@3174.8]
  assign _GEN_81 = _T_637 ? {{1'd0}, _T_1480} : _GEN_80; // @[csr.scala 387:29:Sodor3Stage.fir@3172.6]
  assign _T_1482 = _T_287[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@3179.8]
  assign _T_1483 = {_T_1336,_T_1482}; // @[Cat.scala 30:58:Sodor3Stage.fir@3180.8]
  assign _GEN_82 = _T_643 ? {{1'd0}, _T_1483} : _T_288; // @[csr.scala 386:29:Sodor3Stage.fir@3177.6]
  assign _T_1484 = _T_287[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@3184.8]
  assign _T_1485 = {_T_1484,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@3185.8]
  assign _GEN_83 = _T_641 ? {{1'd0}, _T_1485} : _GEN_82; // @[csr.scala 387:29:Sodor3Stage.fir@3183.6]
  assign _T_1487 = _T_290[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@3190.8]
  assign _T_1488 = {_T_1336,_T_1487}; // @[Cat.scala 30:58:Sodor3Stage.fir@3191.8]
  assign _GEN_84 = _T_647 ? {{1'd0}, _T_1488} : _T_291; // @[csr.scala 386:29:Sodor3Stage.fir@3188.6]
  assign _T_1489 = _T_290[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@3195.8]
  assign _T_1490 = {_T_1489,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@3196.8]
  assign _GEN_85 = _T_645 ? {{1'd0}, _T_1490} : _GEN_84; // @[csr.scala 387:29:Sodor3Stage.fir@3194.6]
  assign _T_1492 = _T_293[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@3201.8]
  assign _T_1493 = {_T_1336,_T_1492}; // @[Cat.scala 30:58:Sodor3Stage.fir@3202.8]
  assign _GEN_86 = _T_651 ? {{1'd0}, _T_1493} : _T_294; // @[csr.scala 386:29:Sodor3Stage.fir@3199.6]
  assign _T_1494 = _T_293[39:32]; // @[csr.scala 387:45:Sodor3Stage.fir@3206.8]
  assign _T_1495 = {_T_1494,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@3207.8]
  assign _GEN_87 = _T_649 ? {{1'd0}, _T_1495} : _GEN_86; // @[csr.scala 387:29:Sodor3Stage.fir@3205.6]
  assign _T_1497 = _T_185[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@3212.8]
  assign _T_1498 = {wdata,_T_1497}; // @[Cat.scala 30:58:Sodor3Stage.fir@3213.8]
  assign _T_1499 = _T_1498[63:6]; // @[util.scala 135:28:Sodor3Stage.fir@3215.8]
  assign _GEN_88 = _T_653 ? _T_1498 : {{57'd0}, _T_177}; // @[csr.scala 386:29:Sodor3Stage.fir@3210.6]
  assign _T_1500 = _T_185[63:32]; // @[csr.scala 387:45:Sodor3Stage.fir@3219.8]
  assign _T_1501 = {_T_1500,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@3220.8]
  assign _T_1502 = _T_1501[63:6]; // @[util.scala 135:28:Sodor3Stage.fir@3222.8]
  assign _GEN_90 = _T_487 ? _T_1501 : _GEN_88; // @[csr.scala 387:29:Sodor3Stage.fir@3218.6]
  assign _T_1504 = _T_197[31:0]; // @[csr.scala 386:72:Sodor3Stage.fir@3227.8]
  assign _T_1505 = {wdata,_T_1504}; // @[Cat.scala 30:58:Sodor3Stage.fir@3228.8]
  assign _T_1506 = _T_1505[63:6]; // @[util.scala 135:28:Sodor3Stage.fir@3230.8]
  assign _GEN_92 = _T_655 ? _T_1505 : {{57'd0}, _T_189}; // @[csr.scala 386:29:Sodor3Stage.fir@3225.6]
  assign _T_1507 = _T_197[63:32]; // @[csr.scala 387:45:Sodor3Stage.fir@3234.8]
  assign _T_1508 = {_T_1507,wdata}; // @[Cat.scala 30:58:Sodor3Stage.fir@3235.8]
  assign _T_1509 = _T_1508[63:6]; // @[util.scala 135:28:Sodor3Stage.fir@3237.8]
  assign _GEN_94 = _T_489 ? _T_1508 : _GEN_92; // @[csr.scala 387:29:Sodor3Stage.fir@3233.6]
  assign _T_1512 = wdata >> 2'h2; // @[csr.scala 368:78:Sodor3Stage.fir@3248.8]
  assign _GEN_469 = {{3'd0}, _T_1512}; // @[csr.scala 368:86:Sodor3Stage.fir@3249.8]
  assign _T_1514 = _GEN_469 << 2'h2; // @[csr.scala 368:86:Sodor3Stage.fir@3249.8]
  assign _GEN_98 = _T_509 ? _T_1514 : {{3'd0}, _GEN_4}; // @[csr.scala 368:40:Sodor3Stage.fir@3246.6]
  assign _T_1516 = wdata & 32'h8000001f; // @[csr.scala 370:62:Sodor3Stage.fir@3256.8]
  assign _GEN_110 = wen ? _GEN_25 : _T_201; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_111 = wen ? _GEN_27 : _T_204; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_112 = wen ? _GEN_29 : _T_207; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_113 = wen ? _GEN_31 : _T_210; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_114 = wen ? _GEN_33 : _T_213; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_115 = wen ? _GEN_35 : _T_216; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_116 = wen ? _GEN_37 : _T_219; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_117 = wen ? _GEN_39 : _T_222; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_118 = wen ? _GEN_41 : _T_225; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_119 = wen ? _GEN_43 : _T_228; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_120 = wen ? _GEN_45 : _T_231; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_121 = wen ? _GEN_47 : _T_234; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_122 = wen ? _GEN_49 : _T_237; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_123 = wen ? _GEN_51 : _T_240; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_124 = wen ? _GEN_53 : _T_243; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_125 = wen ? _GEN_55 : _T_246; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_126 = wen ? _GEN_57 : _T_249; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_127 = wen ? _GEN_59 : _T_252; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_128 = wen ? _GEN_61 : _T_255; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_129 = wen ? _GEN_63 : _T_258; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_130 = wen ? _GEN_65 : _T_261; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_131 = wen ? _GEN_67 : _T_264; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_132 = wen ? _GEN_69 : _T_267; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_133 = wen ? _GEN_71 : _T_270; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_134 = wen ? _GEN_73 : _T_273; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_135 = wen ? _GEN_75 : _T_276; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_136 = wen ? _GEN_77 : _T_279; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_137 = wen ? _GEN_79 : _T_282; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_138 = wen ? _GEN_81 : _T_285; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_139 = wen ? _GEN_83 : _T_288; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_140 = wen ? _GEN_85 : _T_291; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_141 = wen ? _GEN_87 : _T_294; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_142 = wen ? _GEN_90 : {{57'd0}, _T_177}; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_144 = wen ? _GEN_94 : {{57'd0}, _T_189}; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign _GEN_148 = wen ? _GEN_98 : {{3'd0}, _GEN_4}; // @[csr.scala 331:14:Sodor3Stage.fir@2690.4]
  assign io_rw_rdata = _T_1241[31:0];
  assign io_eret = _T_962 | insn_ret;
  assign io_status_debug = 1'h0;
  assign io_status_prv = reg_mstatus_prv;
  assign io_status_sd = 1'h0;
  assign io_status_zero1 = 8'h0;
  assign io_status_tsr = 1'h0;
  assign io_status_tw = 1'h0;
  assign io_status_tvm = 1'h0;
  assign io_status_mxr = 1'h0;
  assign io_status_sum = 1'h0;
  assign io_status_mprv = 1'h0;
  assign io_status_xs = 2'h0;
  assign io_status_fs = 2'h0;
  assign io_status_mpp = 2'h3;
  assign io_status_hpp = 2'h0;
  assign io_status_spp = 1'h0;
  assign io_status_mpie = reg_mstatus_mpie;
  assign io_status_hpie = 1'h0;
  assign io_status_spie = 1'h0;
  assign io_status_upie = 1'h0;
  assign io_status_mie = reg_mstatus_mie;
  assign io_status_hie = 1'h0;
  assign io_status_sie = 1'h0;
  assign io_status_uie = 1'h0;
  assign io_evec = insn_break ? 32'h80000004 : _GEN_13;
  assign _GEN_338_0 = cpu_wen & _T_663;
  assign _GEN_224_0 = io_decode_csr == 12'hb1c;
  assign _GEN_218_0 = io_decode_csr == 12'hb19;
  assign _GEN_323_0 = io_decode_csr == 12'h302;
  assign _GEN_302_0 = io_decode_csr == 12'hb1f;
  assign _GEN_239_0 = io_decode_csr == 12'h7b0;
  assign _GEN_317_0 = io_decode_csr == 12'h7b1;
  assign _GEN_385_0 = cpu_wen & _T_663;
  assign _GEN_197_0 = io_decode_csr == 12'hb8e;
  assign _GEN_296_0 = io_decode_csr == 12'hb1c;
  assign _GEN_203_0 = io_decode_csr == 12'hb91;
  assign _GEN_212_0 = io_decode_csr == 12'hb16;
  assign _GEN_320_0 = io_decode_csr == 12'h340;
  assign _GEN_200_0 = io_decode_csr == 12'hb10;
  assign _GEN_388_0 = _T_970 == 1'h0;
  assign _GEN_191_0 = io_decode_csr == 12'hb8b;
  assign _GEN_181_0 = io_decode_csr == 12'hb86;
  assign _GEN_190_1 = io_decode_csr == 12'hb0b;
  assign _GEN_289_0 = io_decode_csr == 12'hb99;
  assign _GEN_299_0 = io_decode_csr == 12'hb9e;
  assign _GEN_311_0 = io_decode_csr == 12'hb00;
  assign _GEN_206_0 = io_decode_csr == 12'hb13;
  assign _GEN_367_0 = cpu_wen & _T_663;
  assign _GEN_175_0 = io_decode_csr == 12'hb83;
  assign _GEN_305_0 = io_decode_csr == 12'hba1;
  assign _GEN_274_0 = io_decode_csr == 12'hb11;
  assign _GEN_373_0 = cpu_wen & _T_663;
  assign _GEN_376_0 = reset;
  assign _GEN_382_0 = reset;
  assign _GEN_370_0 = reset;
  assign _GEN_349_0 = cpu_wen & _T_663;
  assign _GEN_262_0 = io_decode_csr == 12'hb0b;
  assign _GEN_355_0 = cpu_wen & _T_663;
  assign _GEN_277_0 = io_decode_csr == 12'hb93;
  assign _GEN_194_0 = io_decode_csr == 12'hb0d;
  assign _GEN_184_0 = io_decode_csr == 12'hb08;
  assign _GEN_293_0 = io_decode_csr == 12'hb9b;
  assign _GEN_157_0 = io_decode_csr == 12'hb00;
  assign _GEN_361_0 = cpu_wen & _T_663;
  assign _GEN_256_0 = io_decode_csr == 12'hb08;
  assign _GEN_283_0 = io_decode_csr == 12'hb96;
  assign _GEN_163_0 = io_decode_csr == 12'h344;
  assign _GEN_178_0 = io_decode_csr == 12'hb05;
  assign _GEN_11_0 = io_rw_cmd == 3'h3;
  assign _GEN_259_0 = io_decode_csr == 12'hb8a;
  assign _GEN_358_0 = cpu_wen & _T_663;
  assign _GEN_172_0 = io_decode_csr == 12'h7b2;
  assign _GEN_271_0 = io_decode_csr == 12'hb90;
  assign _GEN_265_0 = io_decode_csr == 12'hb8d;
  assign _GEN_280_0 = io_decode_csr == 12'hb14;
  assign _GEN_160_0 = io_decode_csr == 12'h301;
  assign _GEN_343_0 = cpu_wen & _T_663;
  assign _GEN_379_0 = reset;
  assign _GEN_238_0 = io_decode_csr == 12'h7b0;
  assign _GEN_337_0 = cpu_wen & _T_663;
  assign _GEN_364_0 = cpu_wen & _T_663;
  assign _GEN_244_0 = io_decode_csr == 12'h304;
  assign _GEN_166_0 = io_decode_csr == 12'h341;
  assign _GEN_286_0 = io_decode_csr == 12'hb17;
  assign _GEN_151_0 = insn_ret & _T_980;
  assign _GEN_187_0 = io_decode_csr == 12'hb89;
  assign _GEN_319_1 = io_decode_csr == 12'h341;
  assign _GEN_268_0 = io_decode_csr == 12'hb0e;
  assign _GEN_226_1 = io_decode_csr == 12'hb1d;
  assign _GEN_147_1 = insn_ret & _T_975;
  assign _GEN_352_0 = cpu_wen & _T_663;
  assign _GEN_247_1 = io_decode_csr == 12'hb84;
  assign _GEN_325_1 = cpu_wen & _T_663;
  assign _GEN_169_0 = io_decode_csr == 12'hf14;
  assign _GEN_232_1 = io_decode_csr == 12'hb20;
  assign _GEN_331_1 = cpu_wen & _T_663;
  assign _GEN_346_0 = cpu_wen & _T_663;
  assign _GEN_154_0 = system_insn & _T_676;
  assign _GEN_340_0 = cpu_wen & _T_663;
  assign _GEN_253_0 = io_decode_csr == 12'hb87;
  assign _GEN_211_1 = io_decode_csr == 12'hb95;
  assign _GEN_220_1 = io_decode_csr == 12'hb1a;
  assign _GEN_229_1 = io_decode_csr == 12'hb9e;
  assign _GEN_292_1 = io_decode_csr == 12'hb1a;
  assign _GEN_307_1 = io_decode_csr == 12'hba2;
  assign _GEN_193_1 = io_decode_csr == 12'hb8c;
  assign _GEN_313_1 = io_decode_csr == 12'hb82;
  assign _GEN_328_0 = cpu_wen & _T_663;
  assign _GEN_235_0 = io_decode_csr == 12'hba1;
  assign _GEN_3_3 = _T_177[6];
  assign _GEN_250_0 = io_decode_csr == 12'hb05;
  assign _GEN_208_1 = io_decode_csr == 12'hb14;
  assign _GEN_214_1 = io_decode_csr == 12'hb17;
  assign _GEN_241_0 = io_decode_csr == 12'h300;
  assign _GEN_334_0 = cpu_wen & _T_663;
  assign _GEN_217_0 = io_decode_csr == 12'hb98;
  assign _GEN_316_0 = io_decode_csr == 12'hb02;
  assign _GEN_180_1 = io_decode_csr == 12'hb06;
  assign _GEN_384_1 = cpu_wen & _T_663;
  assign _GEN_301_1 = io_decode_csr == 12'hb9f;
  assign _GEN_196_1 = io_decode_csr == 12'hb0e;
  assign _GEN_186_1 = io_decode_csr == 12'hb09;
  assign _GEN_295_1 = io_decode_csr == 12'hb9c;
  assign _GEN_223_0 = io_decode_csr == 12'hb9b;
  assign _GEN_322_0 = io_decode_csr == 12'h343;
  assign _GEN_279_1 = io_decode_csr == 12'hb94;
  assign _GEN_310_1 = io_decode_csr == 12'hb80;
  assign _GEN_285_1 = io_decode_csr == 12'hb97;
  assign _GEN_202_1 = io_decode_csr == 12'hb11;
  assign _GEN_378_1 = reset;
  assign _GEN_351_1 = cpu_wen & _T_663;
  assign _GEN_387_1 = reset;
  assign _GEN_189_1 = io_decode_csr == 12'hb8a;
  assign _GEN_372_1 = cpu_wen & _T_663;
  assign _GEN_267_1 = io_decode_csr == 12'hb8e;
  assign _GEN_174_1 = io_decode_csr == 12'hb03;
  assign _GEN_205_1 = io_decode_csr == 12'hb92;
  assign _GEN_273_1 = io_decode_csr == 12'hb91;
  assign _GEN_168_1 = io_decode_csr == 12'h342;
  assign _GEN_199_1 = io_decode_csr == 12'hb8f;
  assign _GEN_298_1 = io_decode_csr == 12'hb1d;
  assign _GEN_304_1 = io_decode_csr == 12'hb20;
  assign _GEN_366_1 = cpu_wen & _T_663;
  assign _GEN_360_1 = cpu_wen & _T_663;
  assign _GEN_288_1 = io_decode_csr == 12'hb18;
  assign _GEN_375_1 = cpu_wen & _T_663;
  assign _GEN_255_1 = io_decode_csr == 12'hb88;
  assign _GEN_261_1 = io_decode_csr == 12'hb8b;
  assign _GEN_270_1 = io_decode_csr == 12'hb0f;
  assign _GEN_150_1 = insn_ret & _T_980;
  assign _GEN_333_1 = cpu_wen & _T_663;
  assign _GEN_177_1 = io_decode_csr == 12'hb84;
  assign _GEN_381_1 = reset;
  assign _GEN_276_1 = io_decode_csr == 12'hb12;
  assign _GEN_354_1 = cpu_wen & _T_663;
  assign _GEN_348_1 = cpu_wen & _T_663;
  assign _GEN_249_1 = io_decode_csr == 12'hb85;
  assign _GEN_369_1 = reset;
  assign _GEN_183_1 = io_decode_csr == 12'hb87;
  assign _GEN_282_1 = io_decode_csr == 12'hb15;
  assign _GEN_162_1 = io_decode_csr == 12'h305;
  assign _GEN_156_1 = system_insn & _T_677;
  assign _GEN_165_1 = io_decode_csr == 12'h340;
  assign _GEN_342_1 = cpu_wen & _T_663;
  assign _GEN_264_1 = io_decode_csr == 12'hb0c;
  assign _GEN_159_1 = io_decode_csr == 12'hf13;
  assign _GEN_222_1 = io_decode_csr == 12'hb1b;
  assign _GEN_363_1 = cpu_wen & _T_663;
  assign _GEN_357_1 = cpu_wen & _T_663;
  assign _GEN_321_1 = io_decode_csr == 12'h342;
  assign _GEN_7_3 = _T_664 | _T_665;
  assign _GEN_330_1 = cpu_wen & _T_663;
  assign _GEN_243_1 = io_decode_csr == 12'h304;
  assign _GEN_237_1 = io_decode_csr == 12'hba2;
  assign _GEN_315_1 = io_decode_csr == 12'hb02;
  assign _GEN_336_1 = cpu_wen & _T_663;
  assign _GEN_258_1 = io_decode_csr == 12'hb09;
  assign _GEN_171_1 = io_decode_csr == 12'h7b1;
  assign _GEN_303_1 = io_decode_csr == 12'hba0;
  assign _GEN_146_1 = io_exception;
  assign _GEN_225_1 = io_decode_csr == 12'hb9c;
  assign _GEN_231_1 = io_decode_csr == 12'hb9f;
  assign _GEN_240_1 = io_decode_csr == 12'h300;
  assign _GEN_339_1 = cpu_wen & _T_663;
  assign _GEN_153_1 = insn_ret & _T_980;
  assign _GEN_252_1 = io_decode_csr == 12'hb06;
  assign _GEN_297_1 = io_decode_csr == 12'hb9d;
  assign _GEN_324_1 = cpu_wen & _T_663;
  assign _GEN_219_1 = io_decode_csr == 12'hb99;
  assign _GEN_246_1 = io_decode_csr == 12'hb03;
  assign _GEN_318_1 = io_decode_csr == 12'h7b2;
  assign _GEN_345_1 = cpu_wen & _T_663;
  assign _GEN_204_1 = io_decode_csr == 12'hb12;
  assign _GEN_213_1 = io_decode_csr == 12'hb96;
  assign _GEN_228_1 = io_decode_csr == 12'hb1e;
  assign _GEN_281_1 = io_decode_csr == 12'hb95;
  assign _GEN_234_1 = io_decode_csr == 12'hb21;
  assign _GEN_312_1 = io_decode_csr == 12'hb00;
  assign _GEN_192_1 = io_decode_csr == 12'hb0c;
  assign _GEN_306_1 = io_decode_csr == 12'hb21;
  assign _GEN_207_1 = io_decode_csr == 12'hb93;
  assign _GEN_300_1 = io_decode_csr == 12'hb1e;
  assign _GEN_327_1 = cpu_wen & _T_663;
  assign _GEN_182_1 = io_decode_csr == 12'hb07;
  assign _GEN_291_1 = io_decode_csr == 12'hb9a;
  assign _GEN_290_0 = io_decode_csr == 12'hb19;
  assign _GEN_383_1 = reset;
  assign _GEN_195_1 = io_decode_csr == 12'hb8d;
  assign _GEN_185_1 = io_decode_csr == 12'hb88;
  assign _GEN_179_1 = io_decode_csr == 12'hb85;
  assign _GEN_216_1 = io_decode_csr == 12'hb18;
  assign _GEN_278_1 = io_decode_csr == 12'hb13;
  assign _GEN_201_1 = io_decode_csr == 12'hb90;
  assign _GEN_210_1 = io_decode_csr == 12'hb15;
  assign _GEN_263_1 = io_decode_csr == 12'hb8c;
  assign _GEN_309_1 = io_decode_csr == 12'hb80;
  assign _GEN_164_1 = io_decode_csr == 12'h304;
  assign _GEN_362_1 = cpu_wen & _T_663;
  assign _GEN_377_1 = reset;
  assign _GEN_294_1 = io_decode_csr == 12'hb1b;
  assign _GEN_284_1 = io_decode_csr == 12'hb16;
  assign _GEN_371_1 = reset;
  assign _GEN_260_1 = io_decode_csr == 12'hb0a;
  assign _GEN_266_1 = io_decode_csr == 12'hb0d;
  assign _GEN_380_1 = reset;
  assign _GEN_365_1 = cpu_wen & _T_663;
  assign _GEN_251_1 = io_decode_csr == 12'hb86;
  assign _GEN_15_2 = io_exception;
  assign _GEN_359_1 = cpu_wen & _T_663;
  assign _GEN_152_1 = insn_ret & _T_980;
  assign _GEN_188_1 = io_decode_csr == 12'hb0a;
  assign _GEN_173_1 = io_decode_csr == 12'h302;
  assign _GEN_287_1 = io_decode_csr == 12'hb98;
  assign _GEN_386_1 = reset;
  assign _GEN_245_1 = io_decode_csr == 12'hb83;
  assign _GEN_272_1 = io_decode_csr == 12'hb10;
  assign _GEN_344_1 = cpu_wen & _T_663;
  assign _GEN_198_1 = io_decode_csr == 12'hb0f;
  assign _GEN_167_1 = io_decode_csr == 12'h343;
  assign _GEN_254_1 = io_decode_csr == 12'hb07;
  assign _GEN_161_1 = io_decode_csr == 12'h300;
  assign _GEN_347_1 = cpu_wen & _T_663;
  assign _GEN_170_1 = io_decode_csr == 12'h7b0;
  assign _GEN_275_1 = io_decode_csr == 12'hb92;
  assign _GEN_269_1 = io_decode_csr == 12'hb8f;
  assign _GEN_155_1 = system_insn & _T_676;
  assign _GEN_368_1 = system_insn & _T_677;
  assign _GEN_233_1 = io_decode_csr == 12'hba0;
  assign _GEN_227_1 = io_decode_csr == 12'hb9d;
  assign _GEN_326_1 = cpu_wen & _T_663;
  assign _GEN_149_1 = insn_ret & _T_975;
  assign _GEN_353_1 = cpu_wen & _T_663;
  assign _GEN_248_1 = io_decode_csr == 12'hb04;
  assign _GEN_374_1 = cpu_wen & _T_663;
  assign _GEN_332_1 = cpu_wen & _T_663;
  assign _GEN_176_1 = io_decode_csr == 12'hb04;
  assign _GEN_314_1 = io_decode_csr == 12'hb82;
  assign _GEN_308_1 = io_decode_csr == 12'hb22;
  assign _GEN_341_1 = cpu_wen & _T_663;
  assign _GEN_5_5 = _T_189[6];
  assign _GEN_356_1 = cpu_wen & _T_663;
  assign _GEN_158_1 = io_decode_csr == 12'hb02;
  assign _GEN_209_1 = io_decode_csr == 12'hb94;
  assign _GEN_221_1 = io_decode_csr == 12'hb9a;
  assign _GEN_236_1 = io_decode_csr == 12'hb22;
  assign _GEN_335_1 = cpu_wen & _T_663;
  assign _GEN_329_1 = cpu_wen & _T_663;
  assign _GEN_230_1 = io_decode_csr == 12'hb1f;
  assign _GEN_242_1 = io_decode_csr == 12'h344;
  assign _GEN_257_1 = io_decode_csr == 12'hb89;
  assign _GEN_350_1 = cpu_wen & _T_663;
  assign _GEN_215_1 = io_decode_csr == 12'hb97;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  reg_mstatus_prv = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  reg_mstatus_mpie = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  reg_mstatus_mie = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  reg_mepc = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  reg_mcause = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  reg_mtval = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  reg_mscratch = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  reg_medeleg = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  reg_mip_mtip = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  reg_mip_msip = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  reg_mie_mtip = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  reg_mie_msip = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  _T_176 = _RAND_12[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{$random}};
  _T_180 = _RAND_13[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  _T_188 = _RAND_14[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {2{$random}};
  _T_192 = _RAND_15[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {2{$random}};
  _T_200 = _RAND_16[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {2{$random}};
  _T_203 = _RAND_17[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {2{$random}};
  _T_206 = _RAND_18[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {2{$random}};
  _T_209 = _RAND_19[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {2{$random}};
  _T_212 = _RAND_20[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {2{$random}};
  _T_215 = _RAND_21[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {2{$random}};
  _T_218 = _RAND_22[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {2{$random}};
  _T_221 = _RAND_23[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {2{$random}};
  _T_224 = _RAND_24[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {2{$random}};
  _T_227 = _RAND_25[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {2{$random}};
  _T_230 = _RAND_26[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {2{$random}};
  _T_233 = _RAND_27[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {2{$random}};
  _T_236 = _RAND_28[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {2{$random}};
  _T_239 = _RAND_29[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {2{$random}};
  _T_242 = _RAND_30[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {2{$random}};
  _T_245 = _RAND_31[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {2{$random}};
  _T_248 = _RAND_32[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {2{$random}};
  _T_251 = _RAND_33[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {2{$random}};
  _T_254 = _RAND_34[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {2{$random}};
  _T_257 = _RAND_35[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {2{$random}};
  _T_260 = _RAND_36[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {2{$random}};
  _T_263 = _RAND_37[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {2{$random}};
  _T_266 = _RAND_38[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {2{$random}};
  _T_269 = _RAND_39[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {2{$random}};
  _T_272 = _RAND_40[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {2{$random}};
  _T_275 = _RAND_41[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {2{$random}};
  _T_278 = _RAND_42[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {2{$random}};
  _T_281 = _RAND_43[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {2{$random}};
  _T_284 = _RAND_44[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {2{$random}};
  _T_287 = _RAND_45[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {2{$random}};
  _T_290 = _RAND_46[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {2{$random}};
  _T_293 = _RAND_47[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  reg_dpc = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  reg_dscratch = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  reg_dcsr_ebreakm = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  reg_dcsr_step = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (metaReset) begin
      reg_mstatus_prv <= 2'h0;
    end else begin
      if (reset) begin
        reg_mstatus_prv <= 2'h3;
      end else begin
        if (_T_981) begin
          reg_mstatus_prv <= 2'h3;
        end else begin
          if (_T_976) begin
            reg_mstatus_prv <= 2'h3;
          end
        end
      end
    end
    if (metaReset) begin
      reg_mstatus_mpie <= 1'h0;
    end else begin
      if (reset) begin
        reg_mstatus_mpie <= 1'h0;
      end else begin
        if (wen) begin
          if (_T_499) begin
            reg_mstatus_mpie <= _T_1278;
          end else begin
            if (_T_981) begin
              reg_mstatus_mpie <= 1'h1;
            end
          end
        end else begin
          if (_T_981) begin
            reg_mstatus_mpie <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      reg_mstatus_mie <= 1'h0;
    end else begin
      if (reset) begin
        reg_mstatus_mie <= 1'h0;
      end else begin
        if (wen) begin
          if (_T_499) begin
            reg_mstatus_mie <= _T_1274;
          end else begin
            if (_T_981) begin
              reg_mstatus_mie <= reg_mstatus_mpie;
            end
          end
        end else begin
          if (_T_981) begin
            reg_mstatus_mie <= reg_mstatus_mpie;
          end
        end
      end
    end
    if (metaReset) begin
      reg_mepc <= 32'h0;
    end else begin
      reg_mepc <= _GEN_148[31:0];
    end
    if (metaReset) begin
      reg_mcause <= 32'h0;
    end else begin
      if (wen) begin
        if (_T_513) begin
          reg_mcause <= _T_1516;
        end else begin
          if (insn_break) begin
            reg_mcause <= 32'h3;
          end else begin
            if (insn_call) begin
              reg_mcause <= {{28'd0}, _T_986};
            end else begin
              if (io_exception) begin
                reg_mcause <= 32'h2;
              end
            end
          end
        end
      end else begin
        if (insn_break) begin
          reg_mcause <= 32'h3;
        end else begin
          if (insn_call) begin
            reg_mcause <= {{28'd0}, _T_986};
          end else begin
            if (io_exception) begin
              reg_mcause <= 32'h2;
            end
          end
        end
      end
    end
    if (metaReset) begin
      reg_mtval <= 32'h0;
    end else begin
      if (wen) begin
        if (_T_511) begin
          reg_mtval <= wdata;
        end
      end
    end
    if (metaReset) begin
      reg_mscratch <= 32'h0;
    end else begin
      if (wen) begin
        if (_T_507) begin
          reg_mscratch <= wdata;
        end
      end
    end
    if (metaReset) begin
      reg_medeleg <= 32'h0;
    end else begin
      if (wen) begin
        if (_T_523) begin
          reg_medeleg <= wdata;
        end
      end
    end
    if (metaReset) begin
      reg_mip_mtip <= 1'h0;
    end else begin
      if (reset) begin
        reg_mip_mtip <= 1'h0;
      end else begin
        reg_mip_mtip <= 1'h1;
      end
    end
    if (metaReset) begin
      reg_mip_msip <= 1'h0;
    end else begin
      if (reset) begin
        reg_mip_msip <= 1'h0;
      end else begin
        if (wen) begin
          if (_T_503) begin
            reg_mip_msip <= _T_1302;
          end
        end
      end
    end
    if (metaReset) begin
      reg_mie_mtip <= 1'h0;
    end else begin
      if (reset) begin
        reg_mie_mtip <= 1'h0;
      end else begin
        if (wen) begin
          if (_T_505) begin
            reg_mie_mtip <= _T_1306;
          end
        end
      end
    end
    if (metaReset) begin
      reg_mie_msip <= 1'h0;
    end else begin
      if (reset) begin
        reg_mie_msip <= 1'h0;
      end else begin
        if (wen) begin
          if (_T_505) begin
            reg_mie_msip <= _T_1302;
          end
        end
      end
    end
    if (metaReset) begin
      _T_176 <= 6'h0;
    end else begin
      if (reset) begin
        _T_176 <= 6'h0;
      end else begin
        _T_176 <= _GEN_142[5:0];
      end
    end
    if (metaReset) begin
      _T_180 <= 58'h0;
    end else begin
      if (reset) begin
        _T_180 <= 58'h0;
      end else begin
        if (wen) begin
          if (_T_487) begin
            _T_180 <= _T_1502;
          end else begin
            if (_T_653) begin
              _T_180 <= _T_1499;
            end else begin
              if (_T_181) begin
                _T_180 <= _T_184;
              end
            end
          end
        end else begin
          if (_T_181) begin
            _T_180 <= _T_184;
          end
        end
      end
    end
    if (metaReset) begin
      _T_188 <= 6'h0;
    end else begin
      if (reset) begin
        _T_188 <= 6'h0;
      end else begin
        _T_188 <= _GEN_144[5:0];
      end
    end
    if (metaReset) begin
      _T_192 <= 58'h0;
    end else begin
      if (reset) begin
        _T_192 <= 58'h0;
      end else begin
        if (wen) begin
          if (_T_489) begin
            _T_192 <= _T_1509;
          end else begin
            if (_T_655) begin
              _T_192 <= _T_1506;
            end else begin
              if (_T_193) begin
                _T_192 <= _T_196;
              end
            end
          end
        end else begin
          if (_T_193) begin
            _T_192 <= _T_196;
          end
        end
      end
    end
    if (metaReset) begin
      _T_200 <= 40'h0;
    end else begin
      _T_200 <= _GEN_110[39:0];
    end
    if (metaReset) begin
      _T_203 <= 40'h0;
    end else begin
      _T_203 <= _GEN_111[39:0];
    end
    if (metaReset) begin
      _T_206 <= 40'h0;
    end else begin
      _T_206 <= _GEN_112[39:0];
    end
    if (metaReset) begin
      _T_209 <= 40'h0;
    end else begin
      _T_209 <= _GEN_113[39:0];
    end
    if (metaReset) begin
      _T_212 <= 40'h0;
    end else begin
      _T_212 <= _GEN_114[39:0];
    end
    if (metaReset) begin
      _T_215 <= 40'h0;
    end else begin
      _T_215 <= _GEN_115[39:0];
    end
    if (metaReset) begin
      _T_218 <= 40'h0;
    end else begin
      _T_218 <= _GEN_116[39:0];
    end
    if (metaReset) begin
      _T_221 <= 40'h0;
    end else begin
      _T_221 <= _GEN_117[39:0];
    end
    if (metaReset) begin
      _T_224 <= 40'h0;
    end else begin
      _T_224 <= _GEN_118[39:0];
    end
    if (metaReset) begin
      _T_227 <= 40'h0;
    end else begin
      _T_227 <= _GEN_119[39:0];
    end
    if (metaReset) begin
      _T_230 <= 40'h0;
    end else begin
      _T_230 <= _GEN_120[39:0];
    end
    if (metaReset) begin
      _T_233 <= 40'h0;
    end else begin
      _T_233 <= _GEN_121[39:0];
    end
    if (metaReset) begin
      _T_236 <= 40'h0;
    end else begin
      _T_236 <= _GEN_122[39:0];
    end
    if (metaReset) begin
      _T_239 <= 40'h0;
    end else begin
      _T_239 <= _GEN_123[39:0];
    end
    if (metaReset) begin
      _T_242 <= 40'h0;
    end else begin
      _T_242 <= _GEN_124[39:0];
    end
    if (metaReset) begin
      _T_245 <= 40'h0;
    end else begin
      _T_245 <= _GEN_125[39:0];
    end
    if (metaReset) begin
      _T_248 <= 40'h0;
    end else begin
      _T_248 <= _GEN_126[39:0];
    end
    if (metaReset) begin
      _T_251 <= 40'h0;
    end else begin
      _T_251 <= _GEN_127[39:0];
    end
    if (metaReset) begin
      _T_254 <= 40'h0;
    end else begin
      _T_254 <= _GEN_128[39:0];
    end
    if (metaReset) begin
      _T_257 <= 40'h0;
    end else begin
      _T_257 <= _GEN_129[39:0];
    end
    if (metaReset) begin
      _T_260 <= 40'h0;
    end else begin
      _T_260 <= _GEN_130[39:0];
    end
    if (metaReset) begin
      _T_263 <= 40'h0;
    end else begin
      _T_263 <= _GEN_131[39:0];
    end
    if (metaReset) begin
      _T_266 <= 40'h0;
    end else begin
      _T_266 <= _GEN_132[39:0];
    end
    if (metaReset) begin
      _T_269 <= 40'h0;
    end else begin
      _T_269 <= _GEN_133[39:0];
    end
    if (metaReset) begin
      _T_272 <= 40'h0;
    end else begin
      _T_272 <= _GEN_134[39:0];
    end
    if (metaReset) begin
      _T_275 <= 40'h0;
    end else begin
      _T_275 <= _GEN_135[39:0];
    end
    if (metaReset) begin
      _T_278 <= 40'h0;
    end else begin
      _T_278 <= _GEN_136[39:0];
    end
    if (metaReset) begin
      _T_281 <= 40'h0;
    end else begin
      _T_281 <= _GEN_137[39:0];
    end
    if (metaReset) begin
      _T_284 <= 40'h0;
    end else begin
      _T_284 <= _GEN_138[39:0];
    end
    if (metaReset) begin
      _T_287 <= 40'h0;
    end else begin
      _T_287 <= _GEN_139[39:0];
    end
    if (metaReset) begin
      _T_290 <= 40'h0;
    end else begin
      _T_290 <= _GEN_140[39:0];
    end
    if (metaReset) begin
      _T_293 <= 40'h0;
    end else begin
      _T_293 <= _GEN_141[39:0];
    end
    if (metaReset) begin
      reg_dpc <= 32'h0;
    end else begin
      if (wen) begin
        if (_T_519) begin
          reg_dpc <= wdata;
        end
      end
    end
    if (metaReset) begin
      reg_dscratch <= 32'h0;
    end else begin
      if (wen) begin
        if (_T_521) begin
          reg_dscratch <= wdata;
        end
      end
    end
    if (metaReset) begin
      reg_dcsr_ebreakm <= 1'h0;
    end else begin
      if (reset) begin
        reg_dcsr_ebreakm <= 1'h0;
      end else begin
        if (wen) begin
          if (_T_517) begin
            reg_dcsr_ebreakm <= _T_1262;
          end
        end
      end
    end
    if (metaReset) begin
      reg_dcsr_step <= 1'h0;
    end else begin
      if (reset) begin
        reg_dcsr_step <= 1'h0;
      end else begin
        if (wen) begin
          if (_T_517) begin
            reg_dcsr_step <= _T_1252;
          end
        end
      end
    end
  end
endmodule
module DatPath( // @[:Sodor3Stage.fir@3270.2]
  input         metaReset,
  input         clock, // @[:Sodor3Stage.fir@3271.4]
  input         reset, // @[:Sodor3Stage.fir@3272.4]
  output [31:0] io_imem_req_bits_pc, // @[:Sodor3Stage.fir@3273.4]
  output        io_imem_resp_ready, // @[:Sodor3Stage.fir@3273.4]
  input         io_imem_resp_valid, // @[:Sodor3Stage.fir@3273.4]
  input  [31:0] io_imem_resp_bits_pc, // @[:Sodor3Stage.fir@3273.4]
  input  [31:0] io_imem_resp_bits_inst, // @[:Sodor3Stage.fir@3273.4]
  output [31:0] io_dmem_req_bits_addr, // @[:Sodor3Stage.fir@3273.4]
  output [31:0] io_dmem_req_bits_data, // @[:Sodor3Stage.fir@3273.4]
  output        io_dmem_req_bits_fcn, // @[:Sodor3Stage.fir@3273.4]
  output [2:0]  io_dmem_req_bits_typ, // @[:Sodor3Stage.fir@3273.4]
  input  [31:0] io_dmem_resp_bits_data, // @[:Sodor3Stage.fir@3273.4]
  input         io_ctl_exe_kill, // @[:Sodor3Stage.fir@3273.4]
  input  [2:0]  io_ctl_pc_sel, // @[:Sodor3Stage.fir@3273.4]
  input         io_ctl_brjmp_sel, // @[:Sodor3Stage.fir@3273.4]
  input  [1:0]  io_ctl_op1_sel, // @[:Sodor3Stage.fir@3273.4]
  input  [1:0]  io_ctl_op2_sel, // @[:Sodor3Stage.fir@3273.4]
  input  [3:0]  io_ctl_alu_fun, // @[:Sodor3Stage.fir@3273.4]
  input  [1:0]  io_ctl_wb_sel, // @[:Sodor3Stage.fir@3273.4]
  input         io_ctl_rf_wen, // @[:Sodor3Stage.fir@3273.4]
  input         io_ctl_bypassable, // @[:Sodor3Stage.fir@3273.4]
  input  [2:0]  io_ctl_csr_cmd, // @[:Sodor3Stage.fir@3273.4]
  input         io_ctl_dmem_fcn, // @[:Sodor3Stage.fir@3273.4]
  input  [2:0]  io_ctl_dmem_typ, // @[:Sodor3Stage.fir@3273.4]
  input         io_ctl_exception, // @[:Sodor3Stage.fir@3273.4]
  output        io_dat_br_eq, // @[:Sodor3Stage.fir@3273.4]
  output        io_dat_br_lt, // @[:Sodor3Stage.fir@3273.4]
  output        io_dat_br_ltu, // @[:Sodor3Stage.fir@3273.4]
  output        io_dat_csr_eret, // @[:Sodor3Stage.fir@3273.4]
  output        _GEN_338,
  output        _GEN_224,
  output        _GEN_218,
  output        _GEN_21_0,
  output        _GEN_323,
  output        _GEN_302,
  output        _GEN_6_0,
  output        _GEN_239,
  output        _GEN_317,
  output        _GEN_385,
  output        _GEN_197,
  output        _GEN_12_0,
  output        _GEN_296,
  output        _GEN_9_1,
  output        _GEN_203,
  output        _GEN_0_0,
  output        _GEN_9_2,
  output        _GEN_212,
  output        _GEN_320,
  output        _GEN_200,
  output        _GEN_388,
  output        _GEN_191,
  output        _GEN_181,
  output        _GEN_190_0,
  output        _GEN_15_0,
  output        _GEN_289,
  output        _GEN_299,
  output        _GEN_311,
  output        _GEN_206,
  output        _GEN_367,
  output        _GEN_175,
  output        _GEN_305,
  output        _GEN_274,
  output        _GEN_373,
  output        _GEN_376,
  output        _GEN_382,
  output        _GEN_370,
  output        _GEN_349,
  output        _GEN_262,
  output        _GEN_355,
  output        _GEN_277,
  output        _GEN_194,
  output        _GEN_184,
  output        _GEN_293,
  output        _GEN_157,
  output        _GEN_3_1,
  output        _GEN_361,
  output        _GEN_256,
  output        _GEN_283,
  output        _GEN_163,
  output        _GEN_178,
  output        _GEN_8_0,
  output        _GEN_11_0,
  output        _GEN_259,
  output        _GEN_358,
  output        _GEN_172,
  output        _GEN_271,
  output        _GEN_265,
  output        _GEN_280,
  output        _GEN_160,
  output        _GEN_343,
  output        _GEN_379,
  output        _GEN_238,
  output        _GEN_337,
  output        _GEN_364,
  output        _GEN_244,
  output        _GEN_166,
  output        _GEN_286,
  output        _GEN_151,
  output        _GEN_187,
  output        _GEN_319_0,
  output        _GEN_268,
  output        _GEN_226_0,
  output        _GEN_147_0,
  output        _GEN_352,
  output        _GEN_247_0,
  output        _GEN_325_0,
  output        _GEN_2_0,
  output        _GEN_169,
  output        _GEN_232_0,
  output        _GEN_331_0,
  output        _GEN_346,
  output        _GEN_154,
  output        _GEN_340,
  output        _GEN_253,
  output        _GEN_211_0,
  output        _GEN_220_0,
  output        _GEN_229_0,
  output        _GEN_292_0,
  output        _GEN_307_0,
  output        _GEN_193_0,
  output        _GEN_17_0,
  output        _GEN_11_2,
  output        _GEN_313_0,
  output        _GEN_328,
  output        _GEN_2_1,
  output        _GEN_235,
  output        _GEN_3_3,
  output        _GEN_23_0,
  output        _GEN_250,
  output        _GEN_208_0,
  output        _GEN_214_0,
  output        _GEN_241,
  output        _GEN_5_1,
  output        _GEN_334,
  output        _GEN_217,
  output        _GEN_316,
  output        _GEN_180_0,
  output        _GEN_384_0,
  output        _GEN_301_0,
  output        _GEN_196_0,
  output        _GEN_186_0,
  output        _GEN_295_0,
  output        _GEN_20_0,
  output        _GEN_223,
  output        _GEN_322,
  output        _GEN_5_2,
  output        _GEN_279_0,
  output        _GEN_310_0,
  output        _GEN_285_0,
  output        _GEN_202_0,
  output        _GEN_378_0,
  output        _GEN_351_0,
  output        _GEN_387_0,
  output        _GEN_189_0,
  output        _GEN_14_1,
  output        _GEN_372_0,
  output        _GEN_267_0,
  output        _GEN_174_0,
  output        _GEN_205_0,
  output        _GEN_273_0,
  output        _GEN_168_0,
  output        _GEN_199_0,
  output        _GEN_298_0,
  output        _GEN_304_0,
  output        _GEN_366_0,
  output        _GEN_8_2,
  output        _GEN_360_0,
  output        _GEN_288_0,
  output        _GEN_375_0,
  output        _GEN_255_0,
  output        _GEN_261_0,
  output        _GEN_270_0,
  output        _GEN_150_0,
  output        _GEN_333_0,
  output        _GEN_177_0,
  output        _GEN_381_0,
  output        _GEN_1_2,
  output        _GEN_276_0,
  output        _GEN_10_1,
  output        _GEN_354_0,
  output        _GEN_348_0,
  output        _GEN_249_0,
  output        _GEN_369_0,
  output        _GEN_183_0,
  output        _GEN_282_0,
  output        _GEN_162_0,
  output        _GEN_156_0,
  output        _GEN_165_0,
  output        _GEN_7_2,
  output        _GEN_342_0,
  output        _GEN_264_0,
  output        _GEN_159_0,
  output        _GEN_222_0,
  output        _GEN_363_0,
  output        _GEN_357_0,
  output        _GEN_321_0,
  output        _GEN_7_3,
  output        _GEN_330_0,
  output        _GEN_243_0,
  output        _GEN_237_0,
  output        _GEN_315_0,
  output        _GEN_336_0,
  output        _GEN_258_0,
  output        _GEN_171_0,
  output        _GEN_303_0,
  output        _GEN_146_0,
  output        _GEN_13_1,
  output        _GEN_225_0,
  output        _GEN_7_4,
  output        _GEN_231_0,
  output        _GEN_240_0,
  output        _GEN_339_0,
  output        _GEN_153_0,
  output        _GEN_252_0,
  output        _GEN_297_0,
  output        _GEN_324_0,
  output        _GEN_219_0,
  output        _GEN_1_4,
  output        _GEN_246_0,
  output        _GEN_318_0,
  output        _GEN_345_0,
  output        _GEN_204_0,
  output        _GEN_213_0,
  output        _GEN_228_0,
  output        _GEN_281_0,
  output        _GEN_4_2,
  output        _GEN_0_3,
  output        _GEN_234_0,
  output        _GEN_10_3,
  output        _GEN_312_0,
  output        _GEN_192_0,
  output        _GEN_306_0,
  output        _GEN_207_0,
  output        _GEN_16_0,
  output        _GEN_22_0,
  output        _GEN_300_0,
  output        _GEN_327_0,
  output        _GEN_182_0,
  output        _GEN_291_0,
  output        _GEN_290,
  output        _GEN_4_3,
  output        _GEN_383_0,
  output        _GEN_195_0,
  output        _GEN_185_0,
  output        _GEN_179_0,
  output        _GEN_216_0,
  output        _GEN_278_0,
  output        _GEN_201_0,
  output        _GEN_210_0,
  output        _GEN_263_0,
  output        _GEN_309_0,
  output        _GEN_164_0,
  output        _GEN_362_0,
  output        _GEN_19_0,
  output        _GEN_377_0,
  output        _GEN_294_0,
  output        _GEN_284_0,
  output        _GEN_371_0,
  output        _GEN_260_0,
  output        _GEN_266_0,
  output        _GEN_380_0,
  output        _GEN_365_0,
  output        _GEN_251_0,
  output        _GEN_15_2,
  output        _GEN_359_0,
  output        _GEN_152_0,
  output        _GEN_188_0,
  output        _GEN_173_0,
  output        _GEN_287_0,
  output        _GEN_386_0,
  output        _GEN_245_0,
  output        _GEN_272_0,
  output        _GEN_344_0,
  output        _GEN_198_0,
  output        _GEN_167_0,
  output        _GEN_254_0,
  output        _GEN_3_5,
  output        _GEN_161_0,
  output        _GEN_347_0,
  output        _GEN_170_0,
  output        _GEN_275_0,
  output        _GEN_269_0,
  output        _GEN_155_0,
  output        _GEN_368_0,
  output        _GEN_233_0,
  output        _GEN_227_0,
  output        _GEN_326_0,
  output        _GEN_149_0,
  output        _GEN_353_0,
  output        _GEN_248_0,
  output        _GEN_374_0,
  output        _GEN_332_0,
  output        _GEN_176_0,
  output        _GEN_314_0,
  output        _GEN_308_0,
  output        _GEN_341_0,
  output        _GEN_5_5,
  output        _GEN_18_1,
  output        _GEN_356_0,
  output        _GEN_158_0,
  output        _GEN_209_0,
  output        _GEN_221_0,
  output        _GEN_236_0,
  output        _GEN_335_0,
  output        _GEN_329_0,
  output        _GEN_230_0,
  output        _GEN_242_0,
  output        _GEN_257_0,
  output        _GEN_6_5,
  output        _GEN_350_0,
  output        _GEN_215_0
);
  reg  wb_reg_valid; // @[dpath.scala 52:29:Sodor3Stage.fir@3314.4]
  reg [31:0] _RAND_0;
  reg [1:0] wb_reg_ctrl_wb_sel; // @[dpath.scala 53:29:Sodor3Stage.fir@3315.4]
  reg [31:0] _RAND_1;
  reg  wb_reg_ctrl_rf_wen; // @[dpath.scala 53:29:Sodor3Stage.fir@3315.4]
  reg [31:0] _RAND_2;
  reg  wb_reg_ctrl_bypassable; // @[dpath.scala 53:29:Sodor3Stage.fir@3315.4]
  reg [31:0] _RAND_3;
  reg [2:0] wb_reg_ctrl_csr_cmd; // @[dpath.scala 53:29:Sodor3Stage.fir@3315.4]
  reg [31:0] _RAND_4;
  reg [31:0] wb_reg_alu; // @[dpath.scala 54:29:Sodor3Stage.fir@3316.4]
  reg [31:0] _RAND_5;
  reg [11:0] wb_reg_csr_addr; // @[dpath.scala 55:29:Sodor3Stage.fir@3317.4]
  reg [31:0] _RAND_6;
  reg [4:0] wb_reg_wbaddr; // @[dpath.scala 56:29:Sodor3Stage.fir@3318.4]
  reg [31:0] _RAND_7;
  wire  mem_sparse_metaReset; // @[:Sodor3Stage.fir@3348.4]
  wire  mem_sparse_clock; // @[:Sodor3Stage.fir@3348.4]
  wire  mem_sparse_reset; // @[:Sodor3Stage.fir@3348.4]
  wire [4:0] mem_sparse_io_w_1_addr; // @[:Sodor3Stage.fir@3348.4]
  wire  mem_sparse_io_w_1_en; // @[:Sodor3Stage.fir@3348.4]
  wire [31:0] mem_sparse_io_w_1_data; // @[:Sodor3Stage.fir@3348.4]
  wire [4:0] mem_sparse_io_r_1_addr; // @[:Sodor3Stage.fir@3348.4]
  wire [31:0] mem_sparse_io_r_1_data; // @[:Sodor3Stage.fir@3348.4]
  wire [4:0] mem_sparse_io_r_2_addr; // @[:Sodor3Stage.fir@3348.4]
  wire [31:0] mem_sparse_io_r_2_data; // @[:Sodor3Stage.fir@3348.4]
  wire [3:0] alu_io_fn; // @[dpath.scala 167:20:Sodor3Stage.fir@3429.4]
  wire [31:0] alu_io_in2; // @[dpath.scala 167:20:Sodor3Stage.fir@3429.4]
  wire [31:0] alu_io_in1; // @[dpath.scala 167:20:Sodor3Stage.fir@3429.4]
  wire [31:0] alu_io_out; // @[dpath.scala 167:20:Sodor3Stage.fir@3429.4]
  wire [31:0] alu_io_adder_out; // @[dpath.scala 167:20:Sodor3Stage.fir@3429.4]
  wire  alu__GEN_9_1; // @[dpath.scala 167:20:Sodor3Stage.fir@3429.4]
  wire  alu__GEN_0_0; // @[dpath.scala 167:20:Sodor3Stage.fir@3429.4]
  wire  alu__GEN_8_0; // @[dpath.scala 167:20:Sodor3Stage.fir@3429.4]
  wire  alu__GEN_2_0; // @[dpath.scala 167:20:Sodor3Stage.fir@3429.4]
  wire  alu__GEN_5_1; // @[dpath.scala 167:20:Sodor3Stage.fir@3429.4]
  wire  alu__GEN_10_1; // @[dpath.scala 167:20:Sodor3Stage.fir@3429.4]
  wire  alu__GEN_7_2; // @[dpath.scala 167:20:Sodor3Stage.fir@3429.4]
  wire  alu__GEN_1_4; // @[dpath.scala 167:20:Sodor3Stage.fir@3429.4]
  wire  alu__GEN_4_2; // @[dpath.scala 167:20:Sodor3Stage.fir@3429.4]
  wire  alu__GEN_3_5; // @[dpath.scala 167:20:Sodor3Stage.fir@3429.4]
  wire  alu__GEN_6_5; // @[dpath.scala 167:20:Sodor3Stage.fir@3429.4]
  wire  csr_metaReset; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr_clock; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr_reset; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire [2:0] csr_io_rw_cmd; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire [31:0] csr_io_rw_rdata; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire [31:0] csr_io_rw_wdata; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr_io_eret; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire [11:0] csr_io_decode_csr; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr_io_status_debug; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire [1:0] csr_io_status_prv; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr_io_status_sd; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire [7:0] csr_io_status_zero1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr_io_status_tsr; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr_io_status_tw; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr_io_status_tvm; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr_io_status_mxr; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr_io_status_sum; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr_io_status_mprv; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire [1:0] csr_io_status_xs; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire [1:0] csr_io_status_fs; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire [1:0] csr_io_status_mpp; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire [1:0] csr_io_status_hpp; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr_io_status_spp; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr_io_status_mpie; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr_io_status_hpie; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr_io_status_spie; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr_io_status_upie; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr_io_status_mie; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr_io_status_hie; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr_io_status_sie; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr_io_status_uie; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire [31:0] csr_io_evec; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr_io_exception; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr_io_retire; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire [31:0] csr_io_pc; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_338_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_224_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_218_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_323_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_302_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_239_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_317_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_385_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_197_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_296_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_203_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_212_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_320_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_200_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_388_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_191_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_181_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_190_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_289_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_299_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_311_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_206_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_367_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_175_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_305_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_274_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_373_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_376_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_382_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_370_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_349_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_262_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_355_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_277_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_194_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_184_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_293_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_157_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_361_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_256_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_283_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_163_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_178_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_11_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_259_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_358_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_172_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_271_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_265_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_280_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_160_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_343_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_379_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_238_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_337_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_364_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_244_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_166_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_286_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_151_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_187_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_319_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_268_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_226_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_147_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_352_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_247_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_325_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_169_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_232_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_331_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_346_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_154_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_340_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_253_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_211_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_220_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_229_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_292_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_307_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_193_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_313_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_328_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_235_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_3_3; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_250_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_208_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_214_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_241_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_334_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_217_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_316_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_180_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_384_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_301_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_196_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_186_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_295_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_223_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_322_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_279_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_310_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_285_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_202_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_378_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_351_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_387_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_189_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_372_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_267_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_174_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_205_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_273_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_168_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_199_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_298_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_304_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_366_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_360_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_288_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_375_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_255_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_261_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_270_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_150_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_333_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_177_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_381_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_276_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_354_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_348_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_249_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_369_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_183_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_282_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_162_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_156_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_165_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_342_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_264_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_159_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_222_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_363_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_357_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_321_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_7_3; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_330_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_243_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_237_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_315_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_336_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_258_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_171_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_303_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_146_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_225_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_231_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_240_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_339_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_153_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_252_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_297_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_324_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_219_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_246_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_318_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_345_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_204_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_213_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_228_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_281_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_234_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_312_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_192_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_306_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_207_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_300_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_327_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_182_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_291_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_290_0; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_383_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_195_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_185_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_179_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_216_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_278_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_201_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_210_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_263_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_309_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_164_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_362_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_377_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_294_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_284_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_371_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_260_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_266_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_380_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_365_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_251_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_15_2; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_359_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_152_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_188_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_173_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_287_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_386_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_245_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_272_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_344_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_198_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_167_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_254_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_161_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_347_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_170_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_275_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_269_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_155_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_368_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_233_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_227_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_326_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_149_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_353_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_248_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_374_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_332_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_176_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_314_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_308_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_341_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_5_5; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_356_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_158_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_209_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_221_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_236_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_335_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_329_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_230_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_242_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_257_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_350_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  wire  csr__GEN_215_1; // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
  reg  _T_246; // @[dpath.scala 224:27:Sodor3Stage.fir@3590.4]
  reg [31:0] _RAND_8;
  wire [4:0] exe_rs1_addr; // @[dpath.scala 83:31:Sodor3Stage.fir@3330.4]
  wire  _T_129; // @[dpath.scala 105:42:Sodor3Stage.fir@3334.4]
  wire  _T_131; // @[dpath.scala 105:77:Sodor3Stage.fir@3335.4]
  wire  _T_132; // @[dpath.scala 105:60:Sodor3Stage.fir@3336.4]
  wire  _T_133; // @[dpath.scala 105:85:Sodor3Stage.fir@3337.4]
  wire  _T_135; // @[dpath.scala 105:110:Sodor3Stage.fir@3338.4]
  wire  _T_136; // @[dpath.scala 105:107:Sodor3Stage.fir@3339.4]
  wire [4:0] exe_rs2_addr; // @[dpath.scala 84:31:Sodor3Stage.fir@3331.4]
  wire  _T_137; // @[dpath.scala 106:42:Sodor3Stage.fir@3340.4]
  wire  _T_139; // @[dpath.scala 106:77:Sodor3Stage.fir@3341.4]
  wire  _T_140; // @[dpath.scala 106:60:Sodor3Stage.fir@3342.4]
  wire  _T_141; // @[dpath.scala 106:85:Sodor3Stage.fir@3343.4]
  wire  _T_144; // @[dpath.scala 106:107:Sodor3Stage.fir@3345.4]
  wire  wb_hazard_stall; // @[dpath.scala 105:135:Sodor3Stage.fir@3346.4]
  wire  _T_124; // @[dpath.scala 66:26:Sodor3Stage.fir@3323.4]
  wire  _T_125; // @[dpath.scala 69:36:Sodor3Stage.fir@3325.4]
  wire  _T_126; // @[dpath.scala 70:36:Sodor3Stage.fir@3326.4]
  wire [31:0] exe_jump_reg_target; // @[dpath.scala 63:34:Sodor3Stage.fir@3321.4]
  wire  _T_176; // @[dpath.scala 135:28:Sodor3Stage.fir@3381.4]
  wire [7:0] _T_177; // @[dpath.scala 135:42:Sodor3Stage.fir@3382.4]
  wire [8:0] _T_181; // @[Cat.scala 30:58:Sodor3Stage.fir@3386.4]
  wire  _T_178; // @[dpath.scala 135:59:Sodor3Stage.fir@3383.4]
  wire [9:0] _T_179; // @[dpath.scala 135:73:Sodor3Stage.fir@3384.4]
  wire [10:0] _T_180; // @[Cat.scala 30:58:Sodor3Stage.fir@3385.4]
  wire [19:0] imm_j; // @[Cat.scala 30:58:Sodor3Stage.fir@3387.4]
  wire  _T_199; // @[dpath.scala 142:38:Sodor3Stage.fir@3402.4]
  wire [10:0] _T_203; // @[Bitwise.scala 72:12:Sodor3Stage.fir@3404.4]
  wire [30:0] _T_205; // @[Cat.scala 30:58:Sodor3Stage.fir@3405.4]
  wire [31:0] imm_j_sext; // @[Cat.scala 30:58:Sodor3Stage.fir@3406.4]
  wire  _T_165; // @[dpath.scala 133:42:Sodor3Stage.fir@3372.4]
  wire [1:0] _T_169; // @[Cat.scala 30:58:Sodor3Stage.fir@3376.4]
  wire [5:0] _T_166; // @[dpath.scala 133:55:Sodor3Stage.fir@3373.4]
  wire [3:0] _T_167; // @[dpath.scala 133:72:Sodor3Stage.fir@3374.4]
  wire [9:0] _T_168; // @[Cat.scala 30:58:Sodor3Stage.fir@3375.4]
  wire [11:0] imm_b; // @[Cat.scala 30:58:Sodor3Stage.fir@3377.4]
  wire  _T_192; // @[dpath.scala 141:38:Sodor3Stage.fir@3397.4]
  wire [18:0] _T_196; // @[Bitwise.scala 72:12:Sodor3Stage.fir@3399.4]
  wire [30:0] _T_198; // @[Cat.scala 30:58:Sodor3Stage.fir@3400.4]
  wire [31:0] imm_b_sext; // @[Cat.scala 30:58:Sodor3Stage.fir@3401.4]
  wire [31:0] imm_brjmp; // @[dpath.scala 176:23:Sodor3Stage.fir@3435.4]
  wire [32:0] _T_226; // @[dpath.scala 177:31:Sodor3Stage.fir@3436.4]
  wire [31:0] exe_brjmp_target; // @[dpath.scala 177:31:Sodor3Stage.fir@3437.4]
  wire [31:0] _T_127; // @[dpath.scala 70:21:Sodor3Stage.fir@3327.4]
  wire [31:0] exception_target; // @[dpath.scala 64:34:Sodor3Stage.fir@3322.4]
  wire [4:0] exe_wbaddr; // @[dpath.scala 85:31:Sodor3Stage.fir@3332.4]
  wire  _T_151; // @[dpath.scala 121:47:Sodor3Stage.fir@3355.4]
  wire  _T_311; // @[dpath.scala 238:39:Sodor3Stage.fir@3659.4]
  wire  _T_312; // @[dpath.scala 239:39:Sodor3Stage.fir@3660.4]
  wire  _T_313; // @[dpath.scala 240:39:Sodor3Stage.fir@3661.4]
  wire  _T_314; // @[dpath.scala 241:39:Sodor3Stage.fir@3662.4]
  wire [31:0] _T_315; // @[Mux.scala 61:16:Sodor3Stage.fir@3663.4]
  wire [31:0] _T_316; // @[Mux.scala 61:16:Sodor3Stage.fir@3664.4]
  wire [31:0] _T_317; // @[Mux.scala 61:16:Sodor3Stage.fir@3665.4]
  wire [31:0] regfile__T_156_data; // @[:Sodor3Stage.fir@3348.4]
  wire [31:0] rf_rs1_data; // @[dpath.scala 126:25:Sodor3Stage.fir@3363.4]
  wire [31:0] regfile__T_160_data; // @[:Sodor3Stage.fir@3348.4]
  wire [31:0] rf_rs2_data; // @[dpath.scala 127:25:Sodor3Stage.fir@3366.4]
  wire [11:0] imm_i; // @[dpath.scala 131:24:Sodor3Stage.fir@3367.4]
  wire [6:0] _T_162; // @[dpath.scala 132:28:Sodor3Stage.fir@3368.4]
  wire [11:0] imm_s; // @[Cat.scala 30:58:Sodor3Stage.fir@3370.4]
  wire [19:0] _T_170; // @[dpath.scala 134:28:Sodor3Stage.fir@3378.4]
  wire [31:0] imm_u; // @[Cat.scala 30:58:Sodor3Stage.fir@3380.4]
  wire  _T_182; // @[dpath.scala 139:38:Sodor3Stage.fir@3389.4]
  wire [19:0] _T_186; // @[Bitwise.scala 72:12:Sodor3Stage.fir@3391.4]
  wire [31:0] imm_i_sext; // @[Cat.scala 30:58:Sodor3Stage.fir@3392.4]
  wire  _T_187; // @[dpath.scala 140:38:Sodor3Stage.fir@3393.4]
  wire [19:0] _T_191; // @[Bitwise.scala 72:12:Sodor3Stage.fir@3395.4]
  wire [31:0] imm_s_sext; // @[Cat.scala 30:58:Sodor3Stage.fir@3396.4]
  wire  _T_211; // @[dpath.scala 148:109:Sodor3Stage.fir@3411.4]
  wire [31:0] exe_rs1_data; // @[Mux.scala 61:16:Sodor3Stage.fir@3412.4]
  wire  _T_217; // @[dpath.scala 151:109:Sodor3Stage.fir@3417.4]
  wire [31:0] exe_rs2_data; // @[Mux.scala 61:16:Sodor3Stage.fir@3418.4]
  wire  _T_218; // @[dpath.scala 156:41:Sodor3Stage.fir@3419.4]
  wire  _T_219; // @[dpath.scala 157:41:Sodor3Stage.fir@3420.4]
  wire [31:0] _T_220; // @[dpath.scala 157:25:Sodor3Stage.fir@3421.4]
  wire  _T_221; // @[dpath.scala 160:41:Sodor3Stage.fir@3423.4]
  wire  _T_222; // @[dpath.scala 161:41:Sodor3Stage.fir@3424.4]
  wire  _T_223; // @[dpath.scala 162:41:Sodor3Stage.fir@3425.4]
  wire [31:0] _T_224; // @[dpath.scala 162:25:Sodor3Stage.fir@3426.4]
  wire [31:0] _T_225; // @[dpath.scala 161:25:Sodor3Stage.fir@3427.4]
  wire [31:0] _T_229; // @[:Sodor3Stage.fir@3442.4]
  wire [31:0] _T_230; // @[:Sodor3Stage.fir@3443.4]
  wire  _T_235; // @[dpath.scala 191:48:Sodor3Stage.fir@3450.4]
  wire  _T_237; // @[dpath.scala 199:26:Sodor3Stage.fir@3470.4]
  wire  _T_244; // @[dpath.scala 213:30:Sodor3Stage.fir@3482.4]
  wire [32:0] _T_248; // @[dpath.scala 225:31:Sodor3Stage.fir@3593.4]
  wire [32:0] _T_249; // @[dpath.scala 225:31:Sodor3Stage.fir@3594.4]
  SparseMem mem_sparse ( // @[:Sodor3Stage.fir@3348.4]
    .metaReset(mem_sparse_metaReset),
    .clock(mem_sparse_clock),
    .reset(mem_sparse_reset),
    .io_w_1_addr(mem_sparse_io_w_1_addr),
    .io_w_1_en(mem_sparse_io_w_1_en),
    .io_w_1_data(mem_sparse_io_w_1_data),
    .io_r_1_addr(mem_sparse_io_r_1_addr),
    .io_r_1_data(mem_sparse_io_r_1_data),
    .io_r_2_addr(mem_sparse_io_r_2_addr),
    .io_r_2_data(mem_sparse_io_r_2_data)
  );
  ALU alu ( // @[dpath.scala 167:20:Sodor3Stage.fir@3429.4]
    .io_fn(alu_io_fn),
    .io_in2(alu_io_in2),
    .io_in1(alu_io_in1),
    .io_out(alu_io_out),
    .io_adder_out(alu_io_adder_out),
    ._GEN_9_1(alu__GEN_9_1),
    ._GEN_0_0(alu__GEN_0_0),
    ._GEN_8_0(alu__GEN_8_0),
    ._GEN_2_0(alu__GEN_2_0),
    ._GEN_5_1(alu__GEN_5_1),
    ._GEN_10_1(alu__GEN_10_1),
    ._GEN_7_2(alu__GEN_7_2),
    ._GEN_1_4(alu__GEN_1_4),
    ._GEN_4_2(alu__GEN_4_2),
    ._GEN_3_5(alu__GEN_3_5),
    ._GEN_6_5(alu__GEN_6_5)
  );
  CSRFile csr ( // @[dpath.scala 216:20:Sodor3Stage.fir@3484.4]
    .metaReset(csr_metaReset),
    .clock(csr_clock),
    .reset(csr_reset),
    .io_rw_cmd(csr_io_rw_cmd),
    .io_rw_rdata(csr_io_rw_rdata),
    .io_rw_wdata(csr_io_rw_wdata),
    .io_eret(csr_io_eret),
    .io_decode_csr(csr_io_decode_csr),
    .io_status_debug(csr_io_status_debug),
    .io_status_prv(csr_io_status_prv),
    .io_status_sd(csr_io_status_sd),
    .io_status_zero1(csr_io_status_zero1),
    .io_status_tsr(csr_io_status_tsr),
    .io_status_tw(csr_io_status_tw),
    .io_status_tvm(csr_io_status_tvm),
    .io_status_mxr(csr_io_status_mxr),
    .io_status_sum(csr_io_status_sum),
    .io_status_mprv(csr_io_status_mprv),
    .io_status_xs(csr_io_status_xs),
    .io_status_fs(csr_io_status_fs),
    .io_status_mpp(csr_io_status_mpp),
    .io_status_hpp(csr_io_status_hpp),
    .io_status_spp(csr_io_status_spp),
    .io_status_mpie(csr_io_status_mpie),
    .io_status_hpie(csr_io_status_hpie),
    .io_status_spie(csr_io_status_spie),
    .io_status_upie(csr_io_status_upie),
    .io_status_mie(csr_io_status_mie),
    .io_status_hie(csr_io_status_hie),
    .io_status_sie(csr_io_status_sie),
    .io_status_uie(csr_io_status_uie),
    .io_evec(csr_io_evec),
    .io_exception(csr_io_exception),
    .io_retire(csr_io_retire),
    .io_pc(csr_io_pc),
    ._GEN_338_0(csr__GEN_338_0),
    ._GEN_224_0(csr__GEN_224_0),
    ._GEN_218_0(csr__GEN_218_0),
    ._GEN_323_0(csr__GEN_323_0),
    ._GEN_302_0(csr__GEN_302_0),
    ._GEN_239_0(csr__GEN_239_0),
    ._GEN_317_0(csr__GEN_317_0),
    ._GEN_385_0(csr__GEN_385_0),
    ._GEN_197_0(csr__GEN_197_0),
    ._GEN_296_0(csr__GEN_296_0),
    ._GEN_203_0(csr__GEN_203_0),
    ._GEN_212_0(csr__GEN_212_0),
    ._GEN_320_0(csr__GEN_320_0),
    ._GEN_200_0(csr__GEN_200_0),
    ._GEN_388_0(csr__GEN_388_0),
    ._GEN_191_0(csr__GEN_191_0),
    ._GEN_181_0(csr__GEN_181_0),
    ._GEN_190_1(csr__GEN_190_1),
    ._GEN_289_0(csr__GEN_289_0),
    ._GEN_299_0(csr__GEN_299_0),
    ._GEN_311_0(csr__GEN_311_0),
    ._GEN_206_0(csr__GEN_206_0),
    ._GEN_367_0(csr__GEN_367_0),
    ._GEN_175_0(csr__GEN_175_0),
    ._GEN_305_0(csr__GEN_305_0),
    ._GEN_274_0(csr__GEN_274_0),
    ._GEN_373_0(csr__GEN_373_0),
    ._GEN_376_0(csr__GEN_376_0),
    ._GEN_382_0(csr__GEN_382_0),
    ._GEN_370_0(csr__GEN_370_0),
    ._GEN_349_0(csr__GEN_349_0),
    ._GEN_262_0(csr__GEN_262_0),
    ._GEN_355_0(csr__GEN_355_0),
    ._GEN_277_0(csr__GEN_277_0),
    ._GEN_194_0(csr__GEN_194_0),
    ._GEN_184_0(csr__GEN_184_0),
    ._GEN_293_0(csr__GEN_293_0),
    ._GEN_157_0(csr__GEN_157_0),
    ._GEN_361_0(csr__GEN_361_0),
    ._GEN_256_0(csr__GEN_256_0),
    ._GEN_283_0(csr__GEN_283_0),
    ._GEN_163_0(csr__GEN_163_0),
    ._GEN_178_0(csr__GEN_178_0),
    ._GEN_11_0(csr__GEN_11_0),
    ._GEN_259_0(csr__GEN_259_0),
    ._GEN_358_0(csr__GEN_358_0),
    ._GEN_172_0(csr__GEN_172_0),
    ._GEN_271_0(csr__GEN_271_0),
    ._GEN_265_0(csr__GEN_265_0),
    ._GEN_280_0(csr__GEN_280_0),
    ._GEN_160_0(csr__GEN_160_0),
    ._GEN_343_0(csr__GEN_343_0),
    ._GEN_379_0(csr__GEN_379_0),
    ._GEN_238_0(csr__GEN_238_0),
    ._GEN_337_0(csr__GEN_337_0),
    ._GEN_364_0(csr__GEN_364_0),
    ._GEN_244_0(csr__GEN_244_0),
    ._GEN_166_0(csr__GEN_166_0),
    ._GEN_286_0(csr__GEN_286_0),
    ._GEN_151_0(csr__GEN_151_0),
    ._GEN_187_0(csr__GEN_187_0),
    ._GEN_319_1(csr__GEN_319_1),
    ._GEN_268_0(csr__GEN_268_0),
    ._GEN_226_1(csr__GEN_226_1),
    ._GEN_147_1(csr__GEN_147_1),
    ._GEN_352_0(csr__GEN_352_0),
    ._GEN_247_1(csr__GEN_247_1),
    ._GEN_325_1(csr__GEN_325_1),
    ._GEN_169_0(csr__GEN_169_0),
    ._GEN_232_1(csr__GEN_232_1),
    ._GEN_331_1(csr__GEN_331_1),
    ._GEN_346_0(csr__GEN_346_0),
    ._GEN_154_0(csr__GEN_154_0),
    ._GEN_340_0(csr__GEN_340_0),
    ._GEN_253_0(csr__GEN_253_0),
    ._GEN_211_1(csr__GEN_211_1),
    ._GEN_220_1(csr__GEN_220_1),
    ._GEN_229_1(csr__GEN_229_1),
    ._GEN_292_1(csr__GEN_292_1),
    ._GEN_307_1(csr__GEN_307_1),
    ._GEN_193_1(csr__GEN_193_1),
    ._GEN_313_1(csr__GEN_313_1),
    ._GEN_328_0(csr__GEN_328_0),
    ._GEN_235_0(csr__GEN_235_0),
    ._GEN_3_3(csr__GEN_3_3),
    ._GEN_250_0(csr__GEN_250_0),
    ._GEN_208_1(csr__GEN_208_1),
    ._GEN_214_1(csr__GEN_214_1),
    ._GEN_241_0(csr__GEN_241_0),
    ._GEN_334_0(csr__GEN_334_0),
    ._GEN_217_0(csr__GEN_217_0),
    ._GEN_316_0(csr__GEN_316_0),
    ._GEN_180_1(csr__GEN_180_1),
    ._GEN_384_1(csr__GEN_384_1),
    ._GEN_301_1(csr__GEN_301_1),
    ._GEN_196_1(csr__GEN_196_1),
    ._GEN_186_1(csr__GEN_186_1),
    ._GEN_295_1(csr__GEN_295_1),
    ._GEN_223_0(csr__GEN_223_0),
    ._GEN_322_0(csr__GEN_322_0),
    ._GEN_279_1(csr__GEN_279_1),
    ._GEN_310_1(csr__GEN_310_1),
    ._GEN_285_1(csr__GEN_285_1),
    ._GEN_202_1(csr__GEN_202_1),
    ._GEN_378_1(csr__GEN_378_1),
    ._GEN_351_1(csr__GEN_351_1),
    ._GEN_387_1(csr__GEN_387_1),
    ._GEN_189_1(csr__GEN_189_1),
    ._GEN_372_1(csr__GEN_372_1),
    ._GEN_267_1(csr__GEN_267_1),
    ._GEN_174_1(csr__GEN_174_1),
    ._GEN_205_1(csr__GEN_205_1),
    ._GEN_273_1(csr__GEN_273_1),
    ._GEN_168_1(csr__GEN_168_1),
    ._GEN_199_1(csr__GEN_199_1),
    ._GEN_298_1(csr__GEN_298_1),
    ._GEN_304_1(csr__GEN_304_1),
    ._GEN_366_1(csr__GEN_366_1),
    ._GEN_360_1(csr__GEN_360_1),
    ._GEN_288_1(csr__GEN_288_1),
    ._GEN_375_1(csr__GEN_375_1),
    ._GEN_255_1(csr__GEN_255_1),
    ._GEN_261_1(csr__GEN_261_1),
    ._GEN_270_1(csr__GEN_270_1),
    ._GEN_150_1(csr__GEN_150_1),
    ._GEN_333_1(csr__GEN_333_1),
    ._GEN_177_1(csr__GEN_177_1),
    ._GEN_381_1(csr__GEN_381_1),
    ._GEN_276_1(csr__GEN_276_1),
    ._GEN_354_1(csr__GEN_354_1),
    ._GEN_348_1(csr__GEN_348_1),
    ._GEN_249_1(csr__GEN_249_1),
    ._GEN_369_1(csr__GEN_369_1),
    ._GEN_183_1(csr__GEN_183_1),
    ._GEN_282_1(csr__GEN_282_1),
    ._GEN_162_1(csr__GEN_162_1),
    ._GEN_156_1(csr__GEN_156_1),
    ._GEN_165_1(csr__GEN_165_1),
    ._GEN_342_1(csr__GEN_342_1),
    ._GEN_264_1(csr__GEN_264_1),
    ._GEN_159_1(csr__GEN_159_1),
    ._GEN_222_1(csr__GEN_222_1),
    ._GEN_363_1(csr__GEN_363_1),
    ._GEN_357_1(csr__GEN_357_1),
    ._GEN_321_1(csr__GEN_321_1),
    ._GEN_7_3(csr__GEN_7_3),
    ._GEN_330_1(csr__GEN_330_1),
    ._GEN_243_1(csr__GEN_243_1),
    ._GEN_237_1(csr__GEN_237_1),
    ._GEN_315_1(csr__GEN_315_1),
    ._GEN_336_1(csr__GEN_336_1),
    ._GEN_258_1(csr__GEN_258_1),
    ._GEN_171_1(csr__GEN_171_1),
    ._GEN_303_1(csr__GEN_303_1),
    ._GEN_146_1(csr__GEN_146_1),
    ._GEN_225_1(csr__GEN_225_1),
    ._GEN_231_1(csr__GEN_231_1),
    ._GEN_240_1(csr__GEN_240_1),
    ._GEN_339_1(csr__GEN_339_1),
    ._GEN_153_1(csr__GEN_153_1),
    ._GEN_252_1(csr__GEN_252_1),
    ._GEN_297_1(csr__GEN_297_1),
    ._GEN_324_1(csr__GEN_324_1),
    ._GEN_219_1(csr__GEN_219_1),
    ._GEN_246_1(csr__GEN_246_1),
    ._GEN_318_1(csr__GEN_318_1),
    ._GEN_345_1(csr__GEN_345_1),
    ._GEN_204_1(csr__GEN_204_1),
    ._GEN_213_1(csr__GEN_213_1),
    ._GEN_228_1(csr__GEN_228_1),
    ._GEN_281_1(csr__GEN_281_1),
    ._GEN_234_1(csr__GEN_234_1),
    ._GEN_312_1(csr__GEN_312_1),
    ._GEN_192_1(csr__GEN_192_1),
    ._GEN_306_1(csr__GEN_306_1),
    ._GEN_207_1(csr__GEN_207_1),
    ._GEN_300_1(csr__GEN_300_1),
    ._GEN_327_1(csr__GEN_327_1),
    ._GEN_182_1(csr__GEN_182_1),
    ._GEN_291_1(csr__GEN_291_1),
    ._GEN_290_0(csr__GEN_290_0),
    ._GEN_383_1(csr__GEN_383_1),
    ._GEN_195_1(csr__GEN_195_1),
    ._GEN_185_1(csr__GEN_185_1),
    ._GEN_179_1(csr__GEN_179_1),
    ._GEN_216_1(csr__GEN_216_1),
    ._GEN_278_1(csr__GEN_278_1),
    ._GEN_201_1(csr__GEN_201_1),
    ._GEN_210_1(csr__GEN_210_1),
    ._GEN_263_1(csr__GEN_263_1),
    ._GEN_309_1(csr__GEN_309_1),
    ._GEN_164_1(csr__GEN_164_1),
    ._GEN_362_1(csr__GEN_362_1),
    ._GEN_377_1(csr__GEN_377_1),
    ._GEN_294_1(csr__GEN_294_1),
    ._GEN_284_1(csr__GEN_284_1),
    ._GEN_371_1(csr__GEN_371_1),
    ._GEN_260_1(csr__GEN_260_1),
    ._GEN_266_1(csr__GEN_266_1),
    ._GEN_380_1(csr__GEN_380_1),
    ._GEN_365_1(csr__GEN_365_1),
    ._GEN_251_1(csr__GEN_251_1),
    ._GEN_15_2(csr__GEN_15_2),
    ._GEN_359_1(csr__GEN_359_1),
    ._GEN_152_1(csr__GEN_152_1),
    ._GEN_188_1(csr__GEN_188_1),
    ._GEN_173_1(csr__GEN_173_1),
    ._GEN_287_1(csr__GEN_287_1),
    ._GEN_386_1(csr__GEN_386_1),
    ._GEN_245_1(csr__GEN_245_1),
    ._GEN_272_1(csr__GEN_272_1),
    ._GEN_344_1(csr__GEN_344_1),
    ._GEN_198_1(csr__GEN_198_1),
    ._GEN_167_1(csr__GEN_167_1),
    ._GEN_254_1(csr__GEN_254_1),
    ._GEN_161_1(csr__GEN_161_1),
    ._GEN_347_1(csr__GEN_347_1),
    ._GEN_170_1(csr__GEN_170_1),
    ._GEN_275_1(csr__GEN_275_1),
    ._GEN_269_1(csr__GEN_269_1),
    ._GEN_155_1(csr__GEN_155_1),
    ._GEN_368_1(csr__GEN_368_1),
    ._GEN_233_1(csr__GEN_233_1),
    ._GEN_227_1(csr__GEN_227_1),
    ._GEN_326_1(csr__GEN_326_1),
    ._GEN_149_1(csr__GEN_149_1),
    ._GEN_353_1(csr__GEN_353_1),
    ._GEN_248_1(csr__GEN_248_1),
    ._GEN_374_1(csr__GEN_374_1),
    ._GEN_332_1(csr__GEN_332_1),
    ._GEN_176_1(csr__GEN_176_1),
    ._GEN_314_1(csr__GEN_314_1),
    ._GEN_308_1(csr__GEN_308_1),
    ._GEN_341_1(csr__GEN_341_1),
    ._GEN_5_5(csr__GEN_5_5),
    ._GEN_356_1(csr__GEN_356_1),
    ._GEN_158_1(csr__GEN_158_1),
    ._GEN_209_1(csr__GEN_209_1),
    ._GEN_221_1(csr__GEN_221_1),
    ._GEN_236_1(csr__GEN_236_1),
    ._GEN_335_1(csr__GEN_335_1),
    ._GEN_329_1(csr__GEN_329_1),
    ._GEN_230_1(csr__GEN_230_1),
    ._GEN_242_1(csr__GEN_242_1),
    ._GEN_257_1(csr__GEN_257_1),
    ._GEN_350_1(csr__GEN_350_1),
    ._GEN_215_1(csr__GEN_215_1)
  );
  assign mem_sparse_metaReset = metaReset;
  assign csr_metaReset = metaReset;
  assign exe_rs1_addr = io_imem_resp_bits_inst[19:15]; // @[dpath.scala 83:31:Sodor3Stage.fir@3330.4]
  assign _T_129 = wb_reg_wbaddr == exe_rs1_addr; // @[dpath.scala 105:42:Sodor3Stage.fir@3334.4]
  assign _T_131 = exe_rs1_addr != 5'h0; // @[dpath.scala 105:77:Sodor3Stage.fir@3335.4]
  assign _T_132 = _T_129 & _T_131; // @[dpath.scala 105:60:Sodor3Stage.fir@3336.4]
  assign _T_133 = _T_132 & wb_reg_ctrl_rf_wen; // @[dpath.scala 105:85:Sodor3Stage.fir@3337.4]
  assign _T_135 = wb_reg_ctrl_bypassable == 1'h0; // @[dpath.scala 105:110:Sodor3Stage.fir@3338.4]
  assign _T_136 = _T_133 & _T_135; // @[dpath.scala 105:107:Sodor3Stage.fir@3339.4]
  assign exe_rs2_addr = io_imem_resp_bits_inst[24:20]; // @[dpath.scala 84:31:Sodor3Stage.fir@3331.4]
  assign _T_137 = wb_reg_wbaddr == exe_rs2_addr; // @[dpath.scala 106:42:Sodor3Stage.fir@3340.4]
  assign _T_139 = exe_rs2_addr != 5'h0; // @[dpath.scala 106:77:Sodor3Stage.fir@3341.4]
  assign _T_140 = _T_137 & _T_139; // @[dpath.scala 106:60:Sodor3Stage.fir@3342.4]
  assign _T_141 = _T_140 & wb_reg_ctrl_rf_wen; // @[dpath.scala 106:85:Sodor3Stage.fir@3343.4]
  assign _T_144 = _T_141 & _T_135; // @[dpath.scala 106:107:Sodor3Stage.fir@3345.4]
  assign wb_hazard_stall = _T_136 | _T_144; // @[dpath.scala 105:135:Sodor3Stage.fir@3346.4]
  assign _T_124 = wb_hazard_stall == 1'h0; // @[dpath.scala 66:26:Sodor3Stage.fir@3323.4]
  assign _T_125 = io_ctl_pc_sel == 3'h4; // @[dpath.scala 69:36:Sodor3Stage.fir@3325.4]
  assign _T_126 = io_ctl_pc_sel == 3'h3; // @[dpath.scala 70:36:Sodor3Stage.fir@3326.4]
  assign exe_jump_reg_target = alu_io_adder_out; // @[dpath.scala 63:34:Sodor3Stage.fir@3321.4]
  assign _T_176 = io_imem_resp_bits_inst[31]; // @[dpath.scala 135:28:Sodor3Stage.fir@3381.4]
  assign _T_177 = io_imem_resp_bits_inst[19:12]; // @[dpath.scala 135:42:Sodor3Stage.fir@3382.4]
  assign _T_181 = {_T_176,_T_177}; // @[Cat.scala 30:58:Sodor3Stage.fir@3386.4]
  assign _T_178 = io_imem_resp_bits_inst[20]; // @[dpath.scala 135:59:Sodor3Stage.fir@3383.4]
  assign _T_179 = io_imem_resp_bits_inst[30:21]; // @[dpath.scala 135:73:Sodor3Stage.fir@3384.4]
  assign _T_180 = {_T_178,_T_179}; // @[Cat.scala 30:58:Sodor3Stage.fir@3385.4]
  assign imm_j = {_T_181,_T_180}; // @[Cat.scala 30:58:Sodor3Stage.fir@3387.4]
  assign _T_199 = imm_j[19]; // @[dpath.scala 142:38:Sodor3Stage.fir@3402.4]
  assign _T_203 = _T_199 ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12:Sodor3Stage.fir@3404.4]
  assign _T_205 = {_T_203,imm_j}; // @[Cat.scala 30:58:Sodor3Stage.fir@3405.4]
  assign imm_j_sext = {_T_205,1'h0}; // @[Cat.scala 30:58:Sodor3Stage.fir@3406.4]
  assign _T_165 = io_imem_resp_bits_inst[7]; // @[dpath.scala 133:42:Sodor3Stage.fir@3372.4]
  assign _T_169 = {_T_176,_T_165}; // @[Cat.scala 30:58:Sodor3Stage.fir@3376.4]
  assign _T_166 = io_imem_resp_bits_inst[30:25]; // @[dpath.scala 133:55:Sodor3Stage.fir@3373.4]
  assign _T_167 = io_imem_resp_bits_inst[11:8]; // @[dpath.scala 133:72:Sodor3Stage.fir@3374.4]
  assign _T_168 = {_T_166,_T_167}; // @[Cat.scala 30:58:Sodor3Stage.fir@3375.4]
  assign imm_b = {_T_169,_T_168}; // @[Cat.scala 30:58:Sodor3Stage.fir@3377.4]
  assign _T_192 = imm_b[11]; // @[dpath.scala 141:38:Sodor3Stage.fir@3397.4]
  assign _T_196 = _T_192 ? 19'h7ffff : 19'h0; // @[Bitwise.scala 72:12:Sodor3Stage.fir@3399.4]
  assign _T_198 = {_T_196,imm_b}; // @[Cat.scala 30:58:Sodor3Stage.fir@3400.4]
  assign imm_b_sext = {_T_198,1'h0}; // @[Cat.scala 30:58:Sodor3Stage.fir@3401.4]
  assign imm_brjmp = io_ctl_brjmp_sel ? imm_j_sext : imm_b_sext; // @[dpath.scala 176:23:Sodor3Stage.fir@3435.4]
  assign _T_226 = io_imem_resp_bits_pc + imm_brjmp; // @[dpath.scala 177:31:Sodor3Stage.fir@3436.4]
  assign exe_brjmp_target = _T_226[31:0]; // @[dpath.scala 177:31:Sodor3Stage.fir@3437.4]
  assign _T_127 = _T_126 ? exe_jump_reg_target : exe_brjmp_target; // @[dpath.scala 70:21:Sodor3Stage.fir@3327.4]
  assign exception_target = csr_io_evec; // @[dpath.scala 64:34:Sodor3Stage.fir@3322.4]
  assign exe_wbaddr = io_imem_resp_bits_inst[11:7]; // @[dpath.scala 85:31:Sodor3Stage.fir@3332.4]
  assign _T_151 = wb_reg_wbaddr != 5'h0; // @[dpath.scala 121:47:Sodor3Stage.fir@3355.4]
  assign _T_311 = wb_reg_ctrl_wb_sel == 2'h0; // @[dpath.scala 238:39:Sodor3Stage.fir@3659.4]
  assign _T_312 = wb_reg_ctrl_wb_sel == 2'h1; // @[dpath.scala 239:39:Sodor3Stage.fir@3660.4]
  assign _T_313 = wb_reg_ctrl_wb_sel == 2'h2; // @[dpath.scala 240:39:Sodor3Stage.fir@3661.4]
  assign _T_314 = wb_reg_ctrl_wb_sel == 2'h3; // @[dpath.scala 241:39:Sodor3Stage.fir@3662.4]
  assign _T_315 = _T_314 ? csr_io_rw_rdata : wb_reg_alu; // @[Mux.scala 61:16:Sodor3Stage.fir@3663.4]
  assign _T_316 = _T_313 ? io_imem_resp_bits_pc : _T_315; // @[Mux.scala 61:16:Sodor3Stage.fir@3664.4]
  assign _T_317 = _T_312 ? io_dmem_resp_bits_data : _T_316; // @[Mux.scala 61:16:Sodor3Stage.fir@3665.4]
  assign regfile__T_156_data = mem_sparse_io_r_1_data; // @[:Sodor3Stage.fir@3348.4]
  assign rf_rs1_data = _T_131 ? regfile__T_156_data : 32'h0; // @[dpath.scala 126:25:Sodor3Stage.fir@3363.4]
  assign regfile__T_160_data = mem_sparse_io_r_2_data; // @[:Sodor3Stage.fir@3348.4]
  assign rf_rs2_data = _T_139 ? regfile__T_160_data : 32'h0; // @[dpath.scala 127:25:Sodor3Stage.fir@3366.4]
  assign imm_i = io_imem_resp_bits_inst[31:20]; // @[dpath.scala 131:24:Sodor3Stage.fir@3367.4]
  assign _T_162 = io_imem_resp_bits_inst[31:25]; // @[dpath.scala 132:28:Sodor3Stage.fir@3368.4]
  assign imm_s = {_T_162,exe_wbaddr}; // @[Cat.scala 30:58:Sodor3Stage.fir@3370.4]
  assign _T_170 = io_imem_resp_bits_inst[31:12]; // @[dpath.scala 134:28:Sodor3Stage.fir@3378.4]
  assign imm_u = {_T_170,12'h0}; // @[Cat.scala 30:58:Sodor3Stage.fir@3380.4]
  assign _T_182 = imm_i[11]; // @[dpath.scala 139:38:Sodor3Stage.fir@3389.4]
  assign _T_186 = _T_182 ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12:Sodor3Stage.fir@3391.4]
  assign imm_i_sext = {_T_186,imm_i}; // @[Cat.scala 30:58:Sodor3Stage.fir@3392.4]
  assign _T_187 = imm_s[11]; // @[dpath.scala 140:38:Sodor3Stage.fir@3393.4]
  assign _T_191 = _T_187 ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12:Sodor3Stage.fir@3395.4]
  assign imm_s_sext = {_T_191,imm_s}; // @[Cat.scala 30:58:Sodor3Stage.fir@3396.4]
  assign _T_211 = _T_133 & wb_reg_ctrl_bypassable; // @[dpath.scala 148:109:Sodor3Stage.fir@3411.4]
  assign exe_rs1_data = _T_211 ? wb_reg_alu : rf_rs1_data; // @[Mux.scala 61:16:Sodor3Stage.fir@3412.4]
  assign _T_217 = _T_141 & wb_reg_ctrl_bypassable; // @[dpath.scala 151:109:Sodor3Stage.fir@3417.4]
  assign exe_rs2_data = _T_217 ? wb_reg_alu : rf_rs2_data; // @[Mux.scala 61:16:Sodor3Stage.fir@3418.4]
  assign _T_218 = io_ctl_op1_sel == 2'h2; // @[dpath.scala 156:41:Sodor3Stage.fir@3419.4]
  assign _T_219 = io_ctl_op1_sel == 2'h1; // @[dpath.scala 157:41:Sodor3Stage.fir@3420.4]
  assign _T_220 = _T_219 ? imm_u : exe_rs1_data; // @[dpath.scala 157:25:Sodor3Stage.fir@3421.4]
  assign _T_221 = io_ctl_op2_sel == 2'h1; // @[dpath.scala 160:41:Sodor3Stage.fir@3423.4]
  assign _T_222 = io_ctl_op2_sel == 2'h3; // @[dpath.scala 161:41:Sodor3Stage.fir@3424.4]
  assign _T_223 = io_ctl_op2_sel == 2'h2; // @[dpath.scala 162:41:Sodor3Stage.fir@3425.4]
  assign _T_224 = _T_223 ? imm_s_sext : exe_rs2_data; // @[dpath.scala 162:25:Sodor3Stage.fir@3426.4]
  assign _T_225 = _T_222 ? io_imem_resp_bits_pc : _T_224; // @[dpath.scala 161:25:Sodor3Stage.fir@3427.4]
  assign _T_229 = $signed(exe_rs1_data); // @[:Sodor3Stage.fir@3442.4]
  assign _T_230 = $signed(exe_rs2_data); // @[:Sodor3Stage.fir@3443.4]
  assign _T_235 = io_ctl_dmem_fcn & _T_124; // @[dpath.scala 191:48:Sodor3Stage.fir@3450.4]
  assign _T_237 = wb_hazard_stall | io_ctl_exe_kill; // @[dpath.scala 199:26:Sodor3Stage.fir@3470.4]
  assign _T_244 = io_imem_resp_valid & _T_124; // @[dpath.scala 213:30:Sodor3Stage.fir@3482.4]
  assign _T_248 = io_imem_resp_bits_pc - 32'h4; // @[dpath.scala 225:31:Sodor3Stage.fir@3593.4]
  assign _T_249 = $unsigned(_T_248); // @[dpath.scala 225:31:Sodor3Stage.fir@3594.4]
  assign io_imem_req_bits_pc = _T_125 ? exception_target : _T_127;
  assign io_imem_resp_ready = wb_hazard_stall == 1'h0;
  assign io_dmem_req_bits_addr = alu_io_out;
  assign io_dmem_req_bits_data = _T_217 ? wb_reg_alu : rf_rs2_data;
  assign io_dmem_req_bits_fcn = _T_235 & io_imem_resp_valid;
  assign io_dmem_req_bits_typ = io_ctl_dmem_typ;
  assign io_dat_br_eq = exe_rs1_data == exe_rs2_data;
  assign io_dat_br_lt = $signed(_T_229) < $signed(_T_230);
  assign io_dat_br_ltu = exe_rs1_data < exe_rs2_data;
  assign io_dat_csr_eret = csr_io_eret;
  assign _GEN_338 = csr__GEN_338_0;
  assign _GEN_224 = csr__GEN_224_0;
  assign _GEN_218 = csr__GEN_218_0;
  assign _GEN_21_0 = wb_hazard_stall | io_ctl_exe_kill;
  assign _GEN_323 = csr__GEN_323_0;
  assign _GEN_302 = csr__GEN_302_0;
  assign _GEN_6_0 = wb_reg_ctrl_wb_sel == 2'h1;
  assign _GEN_239 = csr__GEN_239_0;
  assign _GEN_317 = csr__GEN_317_0;
  assign _GEN_385 = csr__GEN_385_0;
  assign _GEN_197 = csr__GEN_197_0;
  assign _GEN_12_0 = _T_141 & wb_reg_ctrl_bypassable;
  assign _GEN_296 = csr__GEN_296_0;
  assign _GEN_9_1 = alu__GEN_9_1;
  assign _GEN_203 = csr__GEN_203_0;
  assign _GEN_0_0 = alu__GEN_0_0;
  assign _GEN_9_2 = imm_i[11];
  assign _GEN_212 = csr__GEN_212_0;
  assign _GEN_320 = csr__GEN_320_0;
  assign _GEN_200 = csr__GEN_200_0;
  assign _GEN_388 = csr__GEN_388_0;
  assign _GEN_191 = csr__GEN_191_0;
  assign _GEN_181 = csr__GEN_181_0;
  assign _GEN_190_0 = csr__GEN_190_1;
  assign _GEN_15_0 = io_ctl_op2_sel == 2'h3;
  assign _GEN_289 = csr__GEN_289_0;
  assign _GEN_299 = csr__GEN_299_0;
  assign _GEN_311 = csr__GEN_311_0;
  assign _GEN_206 = csr__GEN_206_0;
  assign _GEN_367 = csr__GEN_367_0;
  assign _GEN_175 = csr__GEN_175_0;
  assign _GEN_305 = csr__GEN_305_0;
  assign _GEN_274 = csr__GEN_274_0;
  assign _GEN_373 = csr__GEN_373_0;
  assign _GEN_376 = csr__GEN_376_0;
  assign _GEN_382 = csr__GEN_382_0;
  assign _GEN_370 = csr__GEN_370_0;
  assign _GEN_349 = csr__GEN_349_0;
  assign _GEN_262 = csr__GEN_262_0;
  assign _GEN_355 = csr__GEN_355_0;
  assign _GEN_277 = csr__GEN_277_0;
  assign _GEN_194 = csr__GEN_194_0;
  assign _GEN_184 = csr__GEN_184_0;
  assign _GEN_293 = csr__GEN_293_0;
  assign _GEN_157 = csr__GEN_157_0;
  assign _GEN_3_1 = io_ctl_pc_sel == 3'h3;
  assign _GEN_361 = csr__GEN_361_0;
  assign _GEN_256 = csr__GEN_256_0;
  assign _GEN_283 = csr__GEN_283_0;
  assign _GEN_163 = csr__GEN_163_0;
  assign _GEN_178 = csr__GEN_178_0;
  assign _GEN_8_0 = alu__GEN_8_0;
  assign _GEN_11_0 = csr__GEN_11_0;
  assign _GEN_259 = csr__GEN_259_0;
  assign _GEN_358 = csr__GEN_358_0;
  assign _GEN_172 = csr__GEN_172_0;
  assign _GEN_271 = csr__GEN_271_0;
  assign _GEN_265 = csr__GEN_265_0;
  assign _GEN_280 = csr__GEN_280_0;
  assign _GEN_160 = csr__GEN_160_0;
  assign _GEN_343 = csr__GEN_343_0;
  assign _GEN_379 = csr__GEN_379_0;
  assign _GEN_238 = csr__GEN_238_0;
  assign _GEN_337 = csr__GEN_337_0;
  assign _GEN_364 = csr__GEN_364_0;
  assign _GEN_244 = csr__GEN_244_0;
  assign _GEN_166 = csr__GEN_166_0;
  assign _GEN_286 = csr__GEN_286_0;
  assign _GEN_151 = csr__GEN_151_0;
  assign _GEN_187 = csr__GEN_187_0;
  assign _GEN_319_0 = csr__GEN_319_1;
  assign _GEN_268 = csr__GEN_268_0;
  assign _GEN_226_0 = csr__GEN_226_1;
  assign _GEN_147_0 = csr__GEN_147_1;
  assign _GEN_352 = csr__GEN_352_0;
  assign _GEN_247_0 = csr__GEN_247_1;
  assign _GEN_325_0 = csr__GEN_325_1;
  assign _GEN_2_0 = alu__GEN_2_0;
  assign _GEN_169 = csr__GEN_169_0;
  assign _GEN_232_0 = csr__GEN_232_1;
  assign _GEN_331_0 = csr__GEN_331_1;
  assign _GEN_346 = csr__GEN_346_0;
  assign _GEN_154 = csr__GEN_154_0;
  assign _GEN_340 = csr__GEN_340_0;
  assign _GEN_253 = csr__GEN_253_0;
  assign _GEN_211_0 = csr__GEN_211_1;
  assign _GEN_220_0 = csr__GEN_220_1;
  assign _GEN_229_0 = csr__GEN_229_1;
  assign _GEN_292_0 = csr__GEN_292_1;
  assign _GEN_307_0 = csr__GEN_307_1;
  assign _GEN_193_0 = csr__GEN_193_1;
  assign _GEN_17_0 = io_ctl_pc_sel == 3'h4;
  assign _GEN_11_2 = _T_133 & wb_reg_ctrl_bypassable;
  assign _GEN_313_0 = csr__GEN_313_1;
  assign _GEN_328 = csr__GEN_328_0;
  assign _GEN_2_1 = io_ctl_brjmp_sel;
  assign _GEN_235 = csr__GEN_235_0;
  assign _GEN_3_3 = csr__GEN_3_3;
  assign _GEN_23_0 = io_ctl_op1_sel == 2'h2;
  assign _GEN_250 = csr__GEN_250_0;
  assign _GEN_208_0 = csr__GEN_208_1;
  assign _GEN_214_0 = csr__GEN_214_1;
  assign _GEN_241 = csr__GEN_241_0;
  assign _GEN_5_1 = alu__GEN_5_1;
  assign _GEN_334 = csr__GEN_334_0;
  assign _GEN_217 = csr__GEN_217_0;
  assign _GEN_316 = csr__GEN_316_0;
  assign _GEN_180_0 = csr__GEN_180_1;
  assign _GEN_384_0 = csr__GEN_384_1;
  assign _GEN_301_0 = csr__GEN_301_1;
  assign _GEN_196_0 = csr__GEN_196_1;
  assign _GEN_186_0 = csr__GEN_186_1;
  assign _GEN_295_0 = csr__GEN_295_1;
  assign _GEN_20_0 = wb_hazard_stall | io_ctl_exe_kill;
  assign _GEN_223 = csr__GEN_223_0;
  assign _GEN_322 = csr__GEN_322_0;
  assign _GEN_5_2 = wb_reg_ctrl_wb_sel == 2'h2;
  assign _GEN_279_0 = csr__GEN_279_1;
  assign _GEN_310_0 = csr__GEN_310_1;
  assign _GEN_285_0 = csr__GEN_285_1;
  assign _GEN_202_0 = csr__GEN_202_1;
  assign _GEN_378_0 = csr__GEN_378_1;
  assign _GEN_351_0 = csr__GEN_351_1;
  assign _GEN_387_0 = csr__GEN_387_1;
  assign _GEN_189_0 = csr__GEN_189_1;
  assign _GEN_14_1 = io_ctl_op2_sel == 2'h2;
  assign _GEN_372_0 = csr__GEN_372_1;
  assign _GEN_267_0 = csr__GEN_267_1;
  assign _GEN_174_0 = csr__GEN_174_1;
  assign _GEN_205_0 = csr__GEN_205_1;
  assign _GEN_273_0 = csr__GEN_273_1;
  assign _GEN_168_0 = csr__GEN_168_1;
  assign _GEN_199_0 = csr__GEN_199_1;
  assign _GEN_298_0 = csr__GEN_298_1;
  assign _GEN_304_0 = csr__GEN_304_1;
  assign _GEN_366_0 = csr__GEN_366_1;
  assign _GEN_8_2 = exe_rs2_addr != 5'h0;
  assign _GEN_360_0 = csr__GEN_360_1;
  assign _GEN_288_0 = csr__GEN_288_1;
  assign _GEN_375_0 = csr__GEN_375_1;
  assign _GEN_255_0 = csr__GEN_255_1;
  assign _GEN_261_0 = csr__GEN_261_1;
  assign _GEN_270_0 = csr__GEN_270_1;
  assign _GEN_150_0 = csr__GEN_150_1;
  assign _GEN_333_0 = csr__GEN_333_1;
  assign _GEN_177_0 = csr__GEN_177_1;
  assign _GEN_381_0 = csr__GEN_381_1;
  assign _GEN_1_2 = imm_b[11];
  assign _GEN_276_0 = csr__GEN_276_1;
  assign _GEN_10_1 = alu__GEN_10_1;
  assign _GEN_354_0 = csr__GEN_354_1;
  assign _GEN_348_0 = csr__GEN_348_1;
  assign _GEN_249_0 = csr__GEN_249_1;
  assign _GEN_369_0 = csr__GEN_369_1;
  assign _GEN_183_0 = csr__GEN_183_1;
  assign _GEN_282_0 = csr__GEN_282_1;
  assign _GEN_162_0 = csr__GEN_162_1;
  assign _GEN_156_0 = csr__GEN_156_1;
  assign _GEN_165_0 = csr__GEN_165_1;
  assign _GEN_7_2 = alu__GEN_7_2;
  assign _GEN_342_0 = csr__GEN_342_1;
  assign _GEN_264_0 = csr__GEN_264_1;
  assign _GEN_159_0 = csr__GEN_159_1;
  assign _GEN_222_0 = csr__GEN_222_1;
  assign _GEN_363_0 = csr__GEN_363_1;
  assign _GEN_357_0 = csr__GEN_357_1;
  assign _GEN_321_0 = csr__GEN_321_1;
  assign _GEN_7_3 = csr__GEN_7_3;
  assign _GEN_330_0 = csr__GEN_330_1;
  assign _GEN_243_0 = csr__GEN_243_1;
  assign _GEN_237_0 = csr__GEN_237_1;
  assign _GEN_315_0 = csr__GEN_315_1;
  assign _GEN_336_0 = csr__GEN_336_1;
  assign _GEN_258_0 = csr__GEN_258_1;
  assign _GEN_171_0 = csr__GEN_171_1;
  assign _GEN_303_0 = csr__GEN_303_1;
  assign _GEN_146_0 = csr__GEN_146_1;
  assign _GEN_13_1 = io_ctl_op1_sel == 2'h1;
  assign _GEN_225_0 = csr__GEN_225_1;
  assign _GEN_7_4 = exe_rs1_addr != 5'h0;
  assign _GEN_231_0 = csr__GEN_231_1;
  assign _GEN_240_0 = csr__GEN_240_1;
  assign _GEN_339_0 = csr__GEN_339_1;
  assign _GEN_153_0 = csr__GEN_153_1;
  assign _GEN_252_0 = csr__GEN_252_1;
  assign _GEN_297_0 = csr__GEN_297_1;
  assign _GEN_324_0 = csr__GEN_324_1;
  assign _GEN_219_0 = csr__GEN_219_1;
  assign _GEN_1_4 = alu__GEN_1_4;
  assign _GEN_246_0 = csr__GEN_246_1;
  assign _GEN_318_0 = csr__GEN_318_1;
  assign _GEN_345_0 = csr__GEN_345_1;
  assign _GEN_204_0 = csr__GEN_204_1;
  assign _GEN_213_0 = csr__GEN_213_1;
  assign _GEN_228_0 = csr__GEN_228_1;
  assign _GEN_281_0 = csr__GEN_281_1;
  assign _GEN_4_2 = alu__GEN_4_2;
  assign _GEN_0_3 = imm_j[19];
  assign _GEN_234_0 = csr__GEN_234_1;
  assign _GEN_10_3 = imm_s[11];
  assign _GEN_312_0 = csr__GEN_312_1;
  assign _GEN_192_0 = csr__GEN_192_1;
  assign _GEN_306_0 = csr__GEN_306_1;
  assign _GEN_207_0 = csr__GEN_207_1;
  assign _GEN_16_0 = wb_reg_ctrl_wb_sel == 2'h0;
  assign _GEN_22_0 = io_ctl_op2_sel == 2'h1;
  assign _GEN_300_0 = csr__GEN_300_1;
  assign _GEN_327_0 = csr__GEN_327_1;
  assign _GEN_182_0 = csr__GEN_182_1;
  assign _GEN_291_0 = csr__GEN_291_1;
  assign _GEN_290 = csr__GEN_290_0;
  assign _GEN_4_3 = wb_reg_ctrl_wb_sel == 2'h3;
  assign _GEN_383_0 = csr__GEN_383_1;
  assign _GEN_195_0 = csr__GEN_195_1;
  assign _GEN_185_0 = csr__GEN_185_1;
  assign _GEN_179_0 = csr__GEN_179_1;
  assign _GEN_216_0 = csr__GEN_216_1;
  assign _GEN_278_0 = csr__GEN_278_1;
  assign _GEN_201_0 = csr__GEN_201_1;
  assign _GEN_210_0 = csr__GEN_210_1;
  assign _GEN_263_0 = csr__GEN_263_1;
  assign _GEN_309_0 = csr__GEN_309_1;
  assign _GEN_164_0 = csr__GEN_164_1;
  assign _GEN_362_0 = csr__GEN_362_1;
  assign _GEN_19_0 = reset;
  assign _GEN_377_0 = csr__GEN_377_1;
  assign _GEN_294_0 = csr__GEN_294_1;
  assign _GEN_284_0 = csr__GEN_284_1;
  assign _GEN_371_0 = csr__GEN_371_1;
  assign _GEN_260_0 = csr__GEN_260_1;
  assign _GEN_266_0 = csr__GEN_266_1;
  assign _GEN_380_0 = csr__GEN_380_1;
  assign _GEN_365_0 = csr__GEN_365_1;
  assign _GEN_251_0 = csr__GEN_251_1;
  assign _GEN_15_2 = csr__GEN_15_2;
  assign _GEN_359_0 = csr__GEN_359_1;
  assign _GEN_152_0 = csr__GEN_152_1;
  assign _GEN_188_0 = csr__GEN_188_1;
  assign _GEN_173_0 = csr__GEN_173_1;
  assign _GEN_287_0 = csr__GEN_287_1;
  assign _GEN_386_0 = csr__GEN_386_1;
  assign _GEN_245_0 = csr__GEN_245_1;
  assign _GEN_272_0 = csr__GEN_272_1;
  assign _GEN_344_0 = csr__GEN_344_1;
  assign _GEN_198_0 = csr__GEN_198_1;
  assign _GEN_167_0 = csr__GEN_167_1;
  assign _GEN_254_0 = csr__GEN_254_1;
  assign _GEN_3_5 = alu__GEN_3_5;
  assign _GEN_161_0 = csr__GEN_161_1;
  assign _GEN_347_0 = csr__GEN_347_1;
  assign _GEN_170_0 = csr__GEN_170_1;
  assign _GEN_275_0 = csr__GEN_275_1;
  assign _GEN_269_0 = csr__GEN_269_1;
  assign _GEN_155_0 = csr__GEN_155_1;
  assign _GEN_368_0 = csr__GEN_368_1;
  assign _GEN_233_0 = csr__GEN_233_1;
  assign _GEN_227_0 = csr__GEN_227_1;
  assign _GEN_326_0 = csr__GEN_326_1;
  assign _GEN_149_0 = csr__GEN_149_1;
  assign _GEN_353_0 = csr__GEN_353_1;
  assign _GEN_248_0 = csr__GEN_248_1;
  assign _GEN_374_0 = csr__GEN_374_1;
  assign _GEN_332_0 = csr__GEN_332_1;
  assign _GEN_176_0 = csr__GEN_176_1;
  assign _GEN_314_0 = csr__GEN_314_1;
  assign _GEN_308_0 = csr__GEN_308_1;
  assign _GEN_341_0 = csr__GEN_341_1;
  assign _GEN_5_5 = csr__GEN_5_5;
  assign _GEN_18_1 = _T_141 & wb_reg_ctrl_bypassable;
  assign _GEN_356_0 = csr__GEN_356_1;
  assign _GEN_158_0 = csr__GEN_158_1;
  assign _GEN_209_0 = csr__GEN_209_1;
  assign _GEN_221_0 = csr__GEN_221_1;
  assign _GEN_236_0 = csr__GEN_236_1;
  assign _GEN_335_0 = csr__GEN_335_1;
  assign _GEN_329_0 = csr__GEN_329_1;
  assign _GEN_230_0 = csr__GEN_230_1;
  assign _GEN_242_0 = csr__GEN_242_1;
  assign _GEN_257_0 = csr__GEN_257_1;
  assign _GEN_6_5 = alu__GEN_6_5;
  assign _GEN_350_0 = csr__GEN_350_1;
  assign _GEN_215_0 = csr__GEN_215_1;
  assign mem_sparse_clock = clock;
  assign mem_sparse_reset = reset;
  assign mem_sparse_io_w_1_addr = wb_reg_wbaddr;
  assign mem_sparse_io_w_1_en = wb_reg_ctrl_rf_wen & _T_151;
  assign mem_sparse_io_w_1_data = _T_311 ? wb_reg_alu : _T_317;
  assign mem_sparse_io_r_1_addr = io_imem_resp_bits_inst[19:15];
  assign mem_sparse_io_r_2_addr = io_imem_resp_bits_inst[24:20];
  assign alu_io_fn = io_ctl_alu_fun;
  assign alu_io_in2 = _T_221 ? imm_i_sext : _T_225;
  assign alu_io_in1 = _T_218 ? {{27'd0}, exe_rs1_addr} : _T_220;
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_rw_cmd = wb_reg_ctrl_csr_cmd;
  assign csr_io_rw_wdata = wb_reg_alu;
  assign csr_io_decode_csr = wb_reg_csr_addr;
  assign csr_io_exception = _T_246;
  assign csr_io_retire = wb_reg_valid;
  assign csr_io_pc = _T_249[31:0];
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  wb_reg_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  wb_reg_ctrl_wb_sel = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  wb_reg_ctrl_rf_wen = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  wb_reg_ctrl_bypassable = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  wb_reg_ctrl_csr_cmd = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  wb_reg_alu = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  wb_reg_csr_addr = _RAND_6[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  wb_reg_wbaddr = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_246 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (metaReset) begin
      wb_reg_valid <= 1'h0;
    end else begin
      if (reset) begin
        wb_reg_valid <= 1'h0;
      end else begin
        wb_reg_valid <= _T_244;
      end
    end
    if (metaReset) begin
      wb_reg_ctrl_wb_sel <= 2'h0;
    end else begin
      wb_reg_ctrl_wb_sel <= io_ctl_wb_sel;
    end
    if (metaReset) begin
      wb_reg_ctrl_rf_wen <= 1'h0;
    end else begin
      if (_T_237) begin
        wb_reg_ctrl_rf_wen <= 1'h0;
      end else begin
        wb_reg_ctrl_rf_wen <= io_ctl_rf_wen;
      end
    end
    if (metaReset) begin
      wb_reg_ctrl_bypassable <= 1'h0;
    end else begin
      wb_reg_ctrl_bypassable <= io_ctl_bypassable;
    end
    if (metaReset) begin
      wb_reg_ctrl_csr_cmd <= 3'h0;
    end else begin
      if (_T_237) begin
        wb_reg_ctrl_csr_cmd <= 3'h0;
      end else begin
        wb_reg_ctrl_csr_cmd <= io_ctl_csr_cmd;
      end
    end
    if (metaReset) begin
      wb_reg_alu <= 32'h0;
    end else begin
      wb_reg_alu <= alu_io_out;
    end
    if (metaReset) begin
      wb_reg_csr_addr <= 12'h0;
    end else begin
      wb_reg_csr_addr <= io_imem_resp_bits_inst[31:20];
    end
    if (metaReset) begin
      wb_reg_wbaddr <= 5'h0;
    end else begin
      wb_reg_wbaddr <= io_imem_resp_bits_inst[11:7];
    end
    if (metaReset) begin
      _T_246 <= 1'h0;
    end else begin
      _T_246 <= io_ctl_exception;
    end
  end
endmodule
module SparseMem(
  input         metaReset,
  input         clock,
  input         reset,
  input  [4:0]  io_w_1_addr,
  input         io_w_1_en,
  input  [31:0] io_w_1_data,
  input  [4:0]  io_r_1_addr,
  output [31:0] io_r_1_data,
  input  [4:0]  io_r_2_addr,
  output [31:0] io_r_2_data
);
  reg [31:0] mem [0:31];
  reg [31:0] _RAND_0;
  wire [31:0] mem__T_959_data;
  wire [4:0] mem__T_959_addr;
  wire [31:0] mem__T_1124_data;
  wire [4:0] mem__T_1124_addr;
  wire [31:0] mem__T_1289_data;
  wire [4:0] mem__T_1289_addr;
  wire [31:0] mem__T_1484_data;
  wire [4:0] mem__T_1484_addr;
  wire  mem__T_1484_mask;
  wire  mem__T_1484_en;
  wire [31:0] mem__T_1670_data;
  wire [4:0] mem__T_1670_addr;
  wire  mem__T_1670_mask;
  wire  mem__T_1670_en;
  wire [4:0] _GEN_393;
  wire [4:0] _GEN_400;
  wire [4:0] _GEN_404;
  reg  addresses_0_valid;
  reg [31:0] _RAND_1;
  reg [4:0] addresses_0_bits;
  reg [31:0] _RAND_2;
  reg  addresses_1_valid;
  reg [31:0] _RAND_3;
  reg [4:0] addresses_1_bits;
  reg [31:0] _RAND_4;
  reg  addresses_2_valid;
  reg [31:0] _RAND_5;
  reg [4:0] addresses_2_bits;
  reg [31:0] _RAND_6;
  reg  addresses_3_valid;
  reg [31:0] _RAND_7;
  reg [4:0] addresses_3_bits;
  reg [31:0] _RAND_8;
  reg  addresses_4_valid;
  reg [31:0] _RAND_9;
  reg [4:0] addresses_4_bits;
  reg [31:0] _RAND_10;
  reg  addresses_5_valid;
  reg [31:0] _RAND_11;
  reg [4:0] addresses_5_bits;
  reg [31:0] _RAND_12;
  reg  addresses_6_valid;
  reg [31:0] _RAND_13;
  reg [4:0] addresses_6_bits;
  reg [31:0] _RAND_14;
  reg  addresses_7_valid;
  reg [31:0] _RAND_15;
  reg [4:0] addresses_7_bits;
  reg [31:0] _RAND_16;
  reg  addresses_8_valid;
  reg [31:0] _RAND_17;
  reg [4:0] addresses_8_bits;
  reg [31:0] _RAND_18;
  reg  addresses_9_valid;
  reg [31:0] _RAND_19;
  reg [4:0] addresses_9_bits;
  reg [31:0] _RAND_20;
  reg  addresses_10_valid;
  reg [31:0] _RAND_21;
  reg [4:0] addresses_10_bits;
  reg [31:0] _RAND_22;
  reg  addresses_11_valid;
  reg [31:0] _RAND_23;
  reg [4:0] addresses_11_bits;
  reg [31:0] _RAND_24;
  reg  addresses_12_valid;
  reg [31:0] _RAND_25;
  reg [4:0] addresses_12_bits;
  reg [31:0] _RAND_26;
  reg  addresses_13_valid;
  reg [31:0] _RAND_27;
  reg [4:0] addresses_13_bits;
  reg [31:0] _RAND_28;
  reg  addresses_14_valid;
  reg [31:0] _RAND_29;
  reg [4:0] addresses_14_bits;
  reg [31:0] _RAND_30;
  reg  addresses_15_valid;
  reg [31:0] _RAND_31;
  reg [4:0] addresses_15_bits;
  reg [31:0] _RAND_32;
  reg  addresses_16_valid;
  reg [31:0] _RAND_33;
  reg [4:0] addresses_16_bits;
  reg [31:0] _RAND_34;
  reg  addresses_17_valid;
  reg [31:0] _RAND_35;
  reg [4:0] addresses_17_bits;
  reg [31:0] _RAND_36;
  reg  addresses_18_valid;
  reg [31:0] _RAND_37;
  reg [4:0] addresses_18_bits;
  reg [31:0] _RAND_38;
  reg  addresses_19_valid;
  reg [31:0] _RAND_39;
  reg [4:0] addresses_19_bits;
  reg [31:0] _RAND_40;
  reg  addresses_20_valid;
  reg [31:0] _RAND_41;
  reg [4:0] addresses_20_bits;
  reg [31:0] _RAND_42;
  reg  addresses_21_valid;
  reg [31:0] _RAND_43;
  reg [4:0] addresses_21_bits;
  reg [31:0] _RAND_44;
  reg  addresses_22_valid;
  reg [31:0] _RAND_45;
  reg [4:0] addresses_22_bits;
  reg [31:0] _RAND_46;
  reg  addresses_23_valid;
  reg [31:0] _RAND_47;
  reg [4:0] addresses_23_bits;
  reg [31:0] _RAND_48;
  reg  addresses_24_valid;
  reg [31:0] _RAND_49;
  reg [4:0] addresses_24_bits;
  reg [31:0] _RAND_50;
  reg  addresses_25_valid;
  reg [31:0] _RAND_51;
  reg [4:0] addresses_25_bits;
  reg [31:0] _RAND_52;
  reg  addresses_26_valid;
  reg [31:0] _RAND_53;
  reg [4:0] addresses_26_bits;
  reg [31:0] _RAND_54;
  reg  addresses_27_valid;
  reg [31:0] _RAND_55;
  reg [4:0] addresses_27_bits;
  reg [31:0] _RAND_56;
  reg  addresses_28_valid;
  reg [31:0] _RAND_57;
  reg [4:0] addresses_28_bits;
  reg [31:0] _RAND_58;
  reg  addresses_29_valid;
  reg [31:0] _RAND_59;
  reg [4:0] addresses_29_bits;
  reg [31:0] _RAND_60;
  reg  addresses_30_valid;
  reg [31:0] _RAND_61;
  reg [4:0] addresses_30_bits;
  reg [31:0] _RAND_62;
  reg  addresses_31_valid;
  reg [31:0] _RAND_63;
  reg [4:0] addresses_31_bits;
  reg [31:0] _RAND_64;
  reg [5:0] nextAddr;
  reg [31:0] _RAND_65;
  wire  _T_799;
  wire  _T_800;
  wire  _T_801;
  wire  _T_802;
  wire  _T_803;
  wire  _T_804;
  wire  _T_805;
  wire  _T_806;
  wire  _T_807;
  wire  _T_808;
  wire  _T_809;
  wire  _T_810;
  wire  _T_811;
  wire  _T_812;
  wire  _T_813;
  wire  _T_814;
  wire  _T_815;
  wire  _T_816;
  wire  _T_817;
  wire  _T_818;
  wire  _T_819;
  wire  _T_820;
  wire  _T_821;
  wire  _T_822;
  wire  _T_823;
  wire  _T_824;
  wire  _T_825;
  wire  _T_826;
  wire  _T_827;
  wire  _T_828;
  wire  _T_829;
  wire  _T_830;
  wire  _T_831;
  wire  _T_832;
  wire  _T_833;
  wire  _T_834;
  wire  _T_835;
  wire  _T_836;
  wire  _T_837;
  wire  _T_838;
  wire  _T_839;
  wire  _T_840;
  wire  _T_841;
  wire  _T_842;
  wire  _T_843;
  wire  _T_844;
  wire  _T_845;
  wire  _T_846;
  wire  _T_847;
  wire  _T_848;
  wire  _T_849;
  wire  _T_850;
  wire  _T_851;
  wire  _T_852;
  wire  _T_853;
  wire  _T_854;
  wire  _T_855;
  wire  _T_856;
  wire  _T_857;
  wire  _T_858;
  wire  _T_859;
  wire  _T_860;
  wire  _T_861;
  wire  _T_862;
  wire [1:0] _T_900;
  wire [1:0] _T_901;
  wire [3:0] _T_902;
  wire [1:0] _T_903;
  wire [1:0] _T_904;
  wire [3:0] _T_905;
  wire [7:0] _T_906;
  wire [1:0] _T_907;
  wire [1:0] _T_908;
  wire [3:0] _T_909;
  wire [1:0] _T_910;
  wire [1:0] _T_911;
  wire [3:0] _T_912;
  wire [7:0] _T_913;
  wire [15:0] _T_914;
  wire [1:0] _T_915;
  wire [1:0] _T_916;
  wire [3:0] _T_917;
  wire [1:0] _T_918;
  wire [1:0] _T_919;
  wire [3:0] _T_920;
  wire [7:0] _T_921;
  wire [1:0] _T_922;
  wire [1:0] _T_923;
  wire [3:0] _T_924;
  wire [1:0] _T_925;
  wire [1:0] _T_926;
  wire [3:0] _T_927;
  wire [7:0] _T_928;
  wire [15:0] _T_929;
  wire [31:0] _T_930;
  wire  _T_932;
  wire [15:0] _T_933;
  wire [15:0] _T_934;
  wire  _T_936;
  wire [15:0] _T_937;
  wire [7:0] _T_938;
  wire [7:0] _T_939;
  wire  _T_941;
  wire [7:0] _T_942;
  wire [3:0] _T_943;
  wire [3:0] _T_944;
  wire  _T_946;
  wire [3:0] _T_947;
  wire [1:0] _T_948;
  wire [1:0] _T_949;
  wire  _T_951;
  wire [1:0] _T_952;
  wire  _T_953;
  wire [1:0] _T_954;
  wire [2:0] _T_955;
  wire [3:0] _T_956;
  wire  _T_964;
  wire  _T_965;
  wire  _T_966;
  wire  _T_967;
  wire  _T_968;
  wire  _T_969;
  wire  _T_970;
  wire  _T_971;
  wire  _T_972;
  wire  _T_973;
  wire  _T_974;
  wire  _T_975;
  wire  _T_976;
  wire  _T_977;
  wire  _T_978;
  wire  _T_979;
  wire  _T_980;
  wire  _T_981;
  wire  _T_982;
  wire  _T_983;
  wire  _T_984;
  wire  _T_985;
  wire  _T_986;
  wire  _T_987;
  wire  _T_988;
  wire  _T_989;
  wire  _T_990;
  wire  _T_991;
  wire  _T_992;
  wire  _T_993;
  wire  _T_994;
  wire  _T_995;
  wire  _T_996;
  wire  _T_997;
  wire  _T_998;
  wire  _T_999;
  wire  _T_1000;
  wire  _T_1001;
  wire  _T_1002;
  wire  _T_1003;
  wire  _T_1004;
  wire  _T_1005;
  wire  _T_1006;
  wire  _T_1007;
  wire  _T_1008;
  wire  _T_1009;
  wire  _T_1010;
  wire  _T_1011;
  wire  _T_1012;
  wire  _T_1013;
  wire  _T_1014;
  wire  _T_1015;
  wire  _T_1016;
  wire  _T_1017;
  wire  _T_1018;
  wire  _T_1019;
  wire  _T_1020;
  wire  _T_1021;
  wire  _T_1022;
  wire  _T_1023;
  wire  _T_1024;
  wire  _T_1025;
  wire  _T_1026;
  wire  _T_1027;
  wire [1:0] _T_1065;
  wire [1:0] _T_1066;
  wire [3:0] _T_1067;
  wire [1:0] _T_1068;
  wire [1:0] _T_1069;
  wire [3:0] _T_1070;
  wire [7:0] _T_1071;
  wire [1:0] _T_1072;
  wire [1:0] _T_1073;
  wire [3:0] _T_1074;
  wire [1:0] _T_1075;
  wire [1:0] _T_1076;
  wire [3:0] _T_1077;
  wire [7:0] _T_1078;
  wire [15:0] _T_1079;
  wire [1:0] _T_1080;
  wire [1:0] _T_1081;
  wire [3:0] _T_1082;
  wire [1:0] _T_1083;
  wire [1:0] _T_1084;
  wire [3:0] _T_1085;
  wire [7:0] _T_1086;
  wire [1:0] _T_1087;
  wire [1:0] _T_1088;
  wire [3:0] _T_1089;
  wire [1:0] _T_1090;
  wire [1:0] _T_1091;
  wire [3:0] _T_1092;
  wire [7:0] _T_1093;
  wire [15:0] _T_1094;
  wire [31:0] _T_1095;
  wire  _T_1097;
  wire [15:0] _T_1098;
  wire [15:0] _T_1099;
  wire  _T_1101;
  wire [15:0] _T_1102;
  wire [7:0] _T_1103;
  wire [7:0] _T_1104;
  wire  _T_1106;
  wire [7:0] _T_1107;
  wire [3:0] _T_1108;
  wire [3:0] _T_1109;
  wire  _T_1111;
  wire [3:0] _T_1112;
  wire [1:0] _T_1113;
  wire [1:0] _T_1114;
  wire  _T_1116;
  wire [1:0] _T_1117;
  wire  _T_1118;
  wire [1:0] _T_1119;
  wire [2:0] _T_1120;
  wire [3:0] _T_1121;
  wire  _T_1129;
  wire  _T_1130;
  wire  _T_1131;
  wire  _T_1132;
  wire  _T_1133;
  wire  _T_1134;
  wire  _T_1135;
  wire  _T_1136;
  wire  _T_1137;
  wire  _T_1138;
  wire  _T_1139;
  wire  _T_1140;
  wire  _T_1141;
  wire  _T_1142;
  wire  _T_1143;
  wire  _T_1144;
  wire  _T_1145;
  wire  _T_1146;
  wire  _T_1147;
  wire  _T_1148;
  wire  _T_1149;
  wire  _T_1150;
  wire  _T_1151;
  wire  _T_1152;
  wire  _T_1153;
  wire  _T_1154;
  wire  _T_1155;
  wire  _T_1156;
  wire  _T_1157;
  wire  _T_1158;
  wire  _T_1159;
  wire  _T_1160;
  wire  _T_1161;
  wire  _T_1162;
  wire  _T_1163;
  wire  _T_1164;
  wire  _T_1165;
  wire  _T_1166;
  wire  _T_1167;
  wire  _T_1168;
  wire  _T_1169;
  wire  _T_1170;
  wire  _T_1171;
  wire  _T_1172;
  wire  _T_1173;
  wire  _T_1174;
  wire  _T_1175;
  wire  _T_1176;
  wire  _T_1177;
  wire  _T_1178;
  wire  _T_1179;
  wire  _T_1180;
  wire  _T_1181;
  wire  _T_1182;
  wire  _T_1183;
  wire  _T_1184;
  wire  _T_1185;
  wire  _T_1186;
  wire  _T_1187;
  wire  _T_1188;
  wire  _T_1189;
  wire  _T_1190;
  wire  _T_1191;
  wire  _T_1192;
  wire [1:0] _T_1230;
  wire [1:0] _T_1231;
  wire [3:0] _T_1232;
  wire [1:0] _T_1233;
  wire [1:0] _T_1234;
  wire [3:0] _T_1235;
  wire [7:0] _T_1236;
  wire [1:0] _T_1237;
  wire [1:0] _T_1238;
  wire [3:0] _T_1239;
  wire [1:0] _T_1240;
  wire [1:0] _T_1241;
  wire [3:0] _T_1242;
  wire [7:0] _T_1243;
  wire [15:0] _T_1244;
  wire [1:0] _T_1245;
  wire [1:0] _T_1246;
  wire [3:0] _T_1247;
  wire [1:0] _T_1248;
  wire [1:0] _T_1249;
  wire [3:0] _T_1250;
  wire [7:0] _T_1251;
  wire [1:0] _T_1252;
  wire [1:0] _T_1253;
  wire [3:0] _T_1254;
  wire [1:0] _T_1255;
  wire [1:0] _T_1256;
  wire [3:0] _T_1257;
  wire [7:0] _T_1258;
  wire [15:0] _T_1259;
  wire [31:0] _T_1260;
  wire  _T_1262;
  wire [15:0] _T_1263;
  wire [15:0] _T_1264;
  wire  _T_1266;
  wire [15:0] _T_1267;
  wire [7:0] _T_1268;
  wire [7:0] _T_1269;
  wire  _T_1271;
  wire [7:0] _T_1272;
  wire [3:0] _T_1273;
  wire [3:0] _T_1274;
  wire  _T_1276;
  wire [3:0] _T_1277;
  wire [1:0] _T_1278;
  wire [1:0] _T_1279;
  wire  _T_1281;
  wire [1:0] _T_1282;
  wire  _T_1283;
  wire [1:0] _T_1284;
  wire [2:0] _T_1285;
  wire [3:0] _T_1286;
  wire [6:0] _T_1297;
  wire [5:0] _T_1298;
  wire  _T_1463;
  wire [5:0] _T_1465;
  wire  _GEN_264;
  wire  _GEN_265;
  wire  _GEN_266;
  wire  _GEN_267;
  wire  _GEN_268;
  wire  _GEN_269;
  wire  _GEN_270;
  wire  _GEN_271;
  wire  _GEN_272;
  wire  _GEN_273;
  wire  _GEN_274;
  wire  _GEN_275;
  wire  _GEN_276;
  wire  _GEN_277;
  wire  _GEN_278;
  wire  _GEN_279;
  wire  _GEN_280;
  wire  _GEN_281;
  wire  _GEN_282;
  wire  _GEN_283;
  wire  _GEN_284;
  wire  _GEN_285;
  wire  _GEN_286;
  wire  _GEN_287;
  wire  _GEN_288;
  wire  _GEN_289;
  wire  _GEN_290;
  wire  _GEN_291;
  wire  _GEN_292;
  wire  _GEN_293;
  wire  _GEN_294;
  wire  _GEN_295;
  wire [5:0] _T_1488;
  wire  _T_1489;
  wire  _T_1490;
  wire  _T_1491;
  wire  _T_1492;
  wire  _T_1493;
  wire  _T_1494;
  wire  _T_1495;
  wire  _T_1496;
  wire  _T_1497;
  wire  _T_1498;
  wire  _T_1499;
  wire  _T_1500;
  wire  _T_1501;
  wire  _T_1502;
  wire  _T_1503;
  wire  _T_1504;
  wire  _T_1505;
  wire  _T_1506;
  wire  _T_1507;
  wire  _T_1508;
  wire  _T_1509;
  wire  _T_1510;
  wire  _T_1511;
  wire  _T_1512;
  wire  _T_1513;
  wire  _T_1514;
  wire  _T_1515;
  wire  _T_1516;
  wire  _T_1517;
  wire  _T_1518;
  wire  _T_1519;
  wire  _T_1520;
  wire  _T_1521;
  wire  _T_1522;
  wire  _T_1523;
  wire  _T_1524;
  wire  _T_1525;
  wire  _T_1526;
  wire  _T_1527;
  wire  _T_1528;
  wire  _T_1529;
  wire  _T_1530;
  wire  _T_1531;
  wire  _T_1532;
  wire  _T_1533;
  wire  _T_1534;
  wire  _T_1535;
  wire  _T_1536;
  wire  _T_1537;
  wire  _T_1538;
  wire  _T_1539;
  wire  _T_1540;
  wire  _T_1541;
  wire  _T_1542;
  wire  _T_1543;
  wire  _T_1544;
  wire  _T_1545;
  wire  _T_1546;
  wire  _T_1547;
  wire  _T_1548;
  wire  _T_1549;
  wire  _T_1550;
  wire  _T_1551;
  wire  _T_1552;
  wire [1:0] _T_1590;
  wire [1:0] _T_1591;
  wire [3:0] _T_1592;
  wire [1:0] _T_1593;
  wire [1:0] _T_1594;
  wire [3:0] _T_1595;
  wire [7:0] _T_1596;
  wire [1:0] _T_1597;
  wire [1:0] _T_1598;
  wire [3:0] _T_1599;
  wire [1:0] _T_1600;
  wire [1:0] _T_1601;
  wire [3:0] _T_1602;
  wire [7:0] _T_1603;
  wire [15:0] _T_1604;
  wire [1:0] _T_1605;
  wire [1:0] _T_1606;
  wire [3:0] _T_1607;
  wire [1:0] _T_1608;
  wire [1:0] _T_1609;
  wire [3:0] _T_1610;
  wire [7:0] _T_1611;
  wire [1:0] _T_1612;
  wire [1:0] _T_1613;
  wire [3:0] _T_1614;
  wire [1:0] _T_1615;
  wire [1:0] _T_1616;
  wire [3:0] _T_1617;
  wire [7:0] _T_1618;
  wire [15:0] _T_1619;
  wire [31:0] _T_1620;
  wire  _T_1622;
  wire [15:0] _T_1623;
  wire [15:0] _T_1624;
  wire  _T_1626;
  wire [15:0] _T_1627;
  wire [7:0] _T_1628;
  wire [7:0] _T_1629;
  wire  _T_1631;
  wire [7:0] _T_1632;
  wire [3:0] _T_1633;
  wire [3:0] _T_1634;
  wire  _T_1636;
  wire [3:0] _T_1637;
  wire [1:0] _T_1638;
  wire [1:0] _T_1639;
  wire  _T_1641;
  wire [1:0] _T_1642;
  wire  _T_1643;
  wire [1:0] _T_1644;
  wire [2:0] _T_1645;
  wire [3:0] _T_1646;
  wire [4:0] _T_1647;
  wire  _T_1649;
  wire  _T_1650;
  wire [5:0] _T_1651;
  wire  _GEN_328;
  wire  _GEN_329;
  wire  _GEN_330;
  wire  _GEN_331;
  wire  _GEN_332;
  wire  _GEN_333;
  wire  _GEN_334;
  wire  _GEN_335;
  wire  _GEN_336;
  wire  _GEN_337;
  wire  _GEN_338;
  wire  _GEN_339;
  wire  _GEN_340;
  wire  _GEN_341;
  wire  _GEN_342;
  wire  _GEN_343;
  wire  _GEN_344;
  wire  _GEN_345;
  wire  _GEN_346;
  wire  _GEN_347;
  wire  _GEN_348;
  wire  _GEN_349;
  wire  _GEN_350;
  wire  _GEN_351;
  wire  _GEN_352;
  wire  _GEN_353;
  wire  _GEN_354;
  wire  _GEN_355;
  wire  _GEN_356;
  wire  _GEN_357;
  wire  _GEN_358;
  wire  _GEN_359;
  wire [6:0] _T_1672;
  wire [5:0] _T_1673;
  wire [5:0] nextAddrUpdate;
  wire  _T_1675;
  wire  _T_1678;
  wire  _T_1680;
  assign mem__T_959_addr = {_T_936,_T_956};
  assign mem__T_959_data = mem[mem__T_959_addr];
  assign mem__T_1124_addr = {_T_1101,_T_1121};
  assign mem__T_1124_data = mem[mem__T_1124_addr];
  assign mem__T_1289_addr = {_T_1266,_T_1286};
  assign mem__T_1289_data = mem[mem__T_1289_addr];
  assign mem__T_1484_data = 32'h0;
  assign mem__T_1484_addr = _T_1465[4:0];
  assign mem__T_1484_mask = 1'h1;
  assign mem__T_1484_en = 1'h1;
  assign mem__T_1670_data = io_w_1_data;
  assign mem__T_1670_addr = _T_1651[4:0];
  assign mem__T_1670_mask = io_w_1_en;
  assign mem__T_1670_en = io_w_1_en;
  assign _GEN_393 = {_T_936,_T_956};
  assign _GEN_400 = _T_1465[4:0];
  assign _GEN_404 = _T_1651[4:0];
  assign _T_799 = addresses_0_bits == 5'h0;
  assign _T_800 = addresses_0_valid & _T_799;
  assign _T_801 = addresses_1_bits == 5'h0;
  assign _T_802 = addresses_1_valid & _T_801;
  assign _T_803 = addresses_2_bits == 5'h0;
  assign _T_804 = addresses_2_valid & _T_803;
  assign _T_805 = addresses_3_bits == 5'h0;
  assign _T_806 = addresses_3_valid & _T_805;
  assign _T_807 = addresses_4_bits == 5'h0;
  assign _T_808 = addresses_4_valid & _T_807;
  assign _T_809 = addresses_5_bits == 5'h0;
  assign _T_810 = addresses_5_valid & _T_809;
  assign _T_811 = addresses_6_bits == 5'h0;
  assign _T_812 = addresses_6_valid & _T_811;
  assign _T_813 = addresses_7_bits == 5'h0;
  assign _T_814 = addresses_7_valid & _T_813;
  assign _T_815 = addresses_8_bits == 5'h0;
  assign _T_816 = addresses_8_valid & _T_815;
  assign _T_817 = addresses_9_bits == 5'h0;
  assign _T_818 = addresses_9_valid & _T_817;
  assign _T_819 = addresses_10_bits == 5'h0;
  assign _T_820 = addresses_10_valid & _T_819;
  assign _T_821 = addresses_11_bits == 5'h0;
  assign _T_822 = addresses_11_valid & _T_821;
  assign _T_823 = addresses_12_bits == 5'h0;
  assign _T_824 = addresses_12_valid & _T_823;
  assign _T_825 = addresses_13_bits == 5'h0;
  assign _T_826 = addresses_13_valid & _T_825;
  assign _T_827 = addresses_14_bits == 5'h0;
  assign _T_828 = addresses_14_valid & _T_827;
  assign _T_829 = addresses_15_bits == 5'h0;
  assign _T_830 = addresses_15_valid & _T_829;
  assign _T_831 = addresses_16_bits == 5'h0;
  assign _T_832 = addresses_16_valid & _T_831;
  assign _T_833 = addresses_17_bits == 5'h0;
  assign _T_834 = addresses_17_valid & _T_833;
  assign _T_835 = addresses_18_bits == 5'h0;
  assign _T_836 = addresses_18_valid & _T_835;
  assign _T_837 = addresses_19_bits == 5'h0;
  assign _T_838 = addresses_19_valid & _T_837;
  assign _T_839 = addresses_20_bits == 5'h0;
  assign _T_840 = addresses_20_valid & _T_839;
  assign _T_841 = addresses_21_bits == 5'h0;
  assign _T_842 = addresses_21_valid & _T_841;
  assign _T_843 = addresses_22_bits == 5'h0;
  assign _T_844 = addresses_22_valid & _T_843;
  assign _T_845 = addresses_23_bits == 5'h0;
  assign _T_846 = addresses_23_valid & _T_845;
  assign _T_847 = addresses_24_bits == 5'h0;
  assign _T_848 = addresses_24_valid & _T_847;
  assign _T_849 = addresses_25_bits == 5'h0;
  assign _T_850 = addresses_25_valid & _T_849;
  assign _T_851 = addresses_26_bits == 5'h0;
  assign _T_852 = addresses_26_valid & _T_851;
  assign _T_853 = addresses_27_bits == 5'h0;
  assign _T_854 = addresses_27_valid & _T_853;
  assign _T_855 = addresses_28_bits == 5'h0;
  assign _T_856 = addresses_28_valid & _T_855;
  assign _T_857 = addresses_29_bits == 5'h0;
  assign _T_858 = addresses_29_valid & _T_857;
  assign _T_859 = addresses_30_bits == 5'h0;
  assign _T_860 = addresses_30_valid & _T_859;
  assign _T_861 = addresses_31_bits == 5'h0;
  assign _T_862 = addresses_31_valid & _T_861;
  assign _T_900 = {_T_802,_T_800};
  assign _T_901 = {_T_806,_T_804};
  assign _T_902 = {_T_901,_T_900};
  assign _T_903 = {_T_810,_T_808};
  assign _T_904 = {_T_814,_T_812};
  assign _T_905 = {_T_904,_T_903};
  assign _T_906 = {_T_905,_T_902};
  assign _T_907 = {_T_818,_T_816};
  assign _T_908 = {_T_822,_T_820};
  assign _T_909 = {_T_908,_T_907};
  assign _T_910 = {_T_826,_T_824};
  assign _T_911 = {_T_830,_T_828};
  assign _T_912 = {_T_911,_T_910};
  assign _T_913 = {_T_912,_T_909};
  assign _T_914 = {_T_913,_T_906};
  assign _T_915 = {_T_834,_T_832};
  assign _T_916 = {_T_838,_T_836};
  assign _T_917 = {_T_916,_T_915};
  assign _T_918 = {_T_842,_T_840};
  assign _T_919 = {_T_846,_T_844};
  assign _T_920 = {_T_919,_T_918};
  assign _T_921 = {_T_920,_T_917};
  assign _T_922 = {_T_850,_T_848};
  assign _T_923 = {_T_854,_T_852};
  assign _T_924 = {_T_923,_T_922};
  assign _T_925 = {_T_858,_T_856};
  assign _T_926 = {_T_862,_T_860};
  assign _T_927 = {_T_926,_T_925};
  assign _T_928 = {_T_927,_T_924};
  assign _T_929 = {_T_928,_T_921};
  assign _T_930 = {_T_929,_T_914};
  assign _T_932 = _T_930 != 32'h0;
  assign _T_933 = _T_930[31:16];
  assign _T_934 = _T_930[15:0];
  assign _T_936 = _T_933 != 16'h0;
  assign _T_937 = _T_933 | _T_934;
  assign _T_938 = _T_937[15:8];
  assign _T_939 = _T_937[7:0];
  assign _T_941 = _T_938 != 8'h0;
  assign _T_942 = _T_938 | _T_939;
  assign _T_943 = _T_942[7:4];
  assign _T_944 = _T_942[3:0];
  assign _T_946 = _T_943 != 4'h0;
  assign _T_947 = _T_943 | _T_944;
  assign _T_948 = _T_947[3:2];
  assign _T_949 = _T_947[1:0];
  assign _T_951 = _T_948 != 2'h0;
  assign _T_952 = _T_948 | _T_949;
  assign _T_953 = _T_952[1];
  assign _T_954 = {_T_951,_T_953};
  assign _T_955 = {_T_946,_T_954};
  assign _T_956 = {_T_941,_T_955};
  assign _T_964 = addresses_0_bits == io_r_1_addr;
  assign _T_965 = addresses_0_valid & _T_964;
  assign _T_966 = addresses_1_bits == io_r_1_addr;
  assign _T_967 = addresses_1_valid & _T_966;
  assign _T_968 = addresses_2_bits == io_r_1_addr;
  assign _T_969 = addresses_2_valid & _T_968;
  assign _T_970 = addresses_3_bits == io_r_1_addr;
  assign _T_971 = addresses_3_valid & _T_970;
  assign _T_972 = addresses_4_bits == io_r_1_addr;
  assign _T_973 = addresses_4_valid & _T_972;
  assign _T_974 = addresses_5_bits == io_r_1_addr;
  assign _T_975 = addresses_5_valid & _T_974;
  assign _T_976 = addresses_6_bits == io_r_1_addr;
  assign _T_977 = addresses_6_valid & _T_976;
  assign _T_978 = addresses_7_bits == io_r_1_addr;
  assign _T_979 = addresses_7_valid & _T_978;
  assign _T_980 = addresses_8_bits == io_r_1_addr;
  assign _T_981 = addresses_8_valid & _T_980;
  assign _T_982 = addresses_9_bits == io_r_1_addr;
  assign _T_983 = addresses_9_valid & _T_982;
  assign _T_984 = addresses_10_bits == io_r_1_addr;
  assign _T_985 = addresses_10_valid & _T_984;
  assign _T_986 = addresses_11_bits == io_r_1_addr;
  assign _T_987 = addresses_11_valid & _T_986;
  assign _T_988 = addresses_12_bits == io_r_1_addr;
  assign _T_989 = addresses_12_valid & _T_988;
  assign _T_990 = addresses_13_bits == io_r_1_addr;
  assign _T_991 = addresses_13_valid & _T_990;
  assign _T_992 = addresses_14_bits == io_r_1_addr;
  assign _T_993 = addresses_14_valid & _T_992;
  assign _T_994 = addresses_15_bits == io_r_1_addr;
  assign _T_995 = addresses_15_valid & _T_994;
  assign _T_996 = addresses_16_bits == io_r_1_addr;
  assign _T_997 = addresses_16_valid & _T_996;
  assign _T_998 = addresses_17_bits == io_r_1_addr;
  assign _T_999 = addresses_17_valid & _T_998;
  assign _T_1000 = addresses_18_bits == io_r_1_addr;
  assign _T_1001 = addresses_18_valid & _T_1000;
  assign _T_1002 = addresses_19_bits == io_r_1_addr;
  assign _T_1003 = addresses_19_valid & _T_1002;
  assign _T_1004 = addresses_20_bits == io_r_1_addr;
  assign _T_1005 = addresses_20_valid & _T_1004;
  assign _T_1006 = addresses_21_bits == io_r_1_addr;
  assign _T_1007 = addresses_21_valid & _T_1006;
  assign _T_1008 = addresses_22_bits == io_r_1_addr;
  assign _T_1009 = addresses_22_valid & _T_1008;
  assign _T_1010 = addresses_23_bits == io_r_1_addr;
  assign _T_1011 = addresses_23_valid & _T_1010;
  assign _T_1012 = addresses_24_bits == io_r_1_addr;
  assign _T_1013 = addresses_24_valid & _T_1012;
  assign _T_1014 = addresses_25_bits == io_r_1_addr;
  assign _T_1015 = addresses_25_valid & _T_1014;
  assign _T_1016 = addresses_26_bits == io_r_1_addr;
  assign _T_1017 = addresses_26_valid & _T_1016;
  assign _T_1018 = addresses_27_bits == io_r_1_addr;
  assign _T_1019 = addresses_27_valid & _T_1018;
  assign _T_1020 = addresses_28_bits == io_r_1_addr;
  assign _T_1021 = addresses_28_valid & _T_1020;
  assign _T_1022 = addresses_29_bits == io_r_1_addr;
  assign _T_1023 = addresses_29_valid & _T_1022;
  assign _T_1024 = addresses_30_bits == io_r_1_addr;
  assign _T_1025 = addresses_30_valid & _T_1024;
  assign _T_1026 = addresses_31_bits == io_r_1_addr;
  assign _T_1027 = addresses_31_valid & _T_1026;
  assign _T_1065 = {_T_967,_T_965};
  assign _T_1066 = {_T_971,_T_969};
  assign _T_1067 = {_T_1066,_T_1065};
  assign _T_1068 = {_T_975,_T_973};
  assign _T_1069 = {_T_979,_T_977};
  assign _T_1070 = {_T_1069,_T_1068};
  assign _T_1071 = {_T_1070,_T_1067};
  assign _T_1072 = {_T_983,_T_981};
  assign _T_1073 = {_T_987,_T_985};
  assign _T_1074 = {_T_1073,_T_1072};
  assign _T_1075 = {_T_991,_T_989};
  assign _T_1076 = {_T_995,_T_993};
  assign _T_1077 = {_T_1076,_T_1075};
  assign _T_1078 = {_T_1077,_T_1074};
  assign _T_1079 = {_T_1078,_T_1071};
  assign _T_1080 = {_T_999,_T_997};
  assign _T_1081 = {_T_1003,_T_1001};
  assign _T_1082 = {_T_1081,_T_1080};
  assign _T_1083 = {_T_1007,_T_1005};
  assign _T_1084 = {_T_1011,_T_1009};
  assign _T_1085 = {_T_1084,_T_1083};
  assign _T_1086 = {_T_1085,_T_1082};
  assign _T_1087 = {_T_1015,_T_1013};
  assign _T_1088 = {_T_1019,_T_1017};
  assign _T_1089 = {_T_1088,_T_1087};
  assign _T_1090 = {_T_1023,_T_1021};
  assign _T_1091 = {_T_1027,_T_1025};
  assign _T_1092 = {_T_1091,_T_1090};
  assign _T_1093 = {_T_1092,_T_1089};
  assign _T_1094 = {_T_1093,_T_1086};
  assign _T_1095 = {_T_1094,_T_1079};
  assign _T_1097 = _T_1095 != 32'h0;
  assign _T_1098 = _T_1095[31:16];
  assign _T_1099 = _T_1095[15:0];
  assign _T_1101 = _T_1098 != 16'h0;
  assign _T_1102 = _T_1098 | _T_1099;
  assign _T_1103 = _T_1102[15:8];
  assign _T_1104 = _T_1102[7:0];
  assign _T_1106 = _T_1103 != 8'h0;
  assign _T_1107 = _T_1103 | _T_1104;
  assign _T_1108 = _T_1107[7:4];
  assign _T_1109 = _T_1107[3:0];
  assign _T_1111 = _T_1108 != 4'h0;
  assign _T_1112 = _T_1108 | _T_1109;
  assign _T_1113 = _T_1112[3:2];
  assign _T_1114 = _T_1112[1:0];
  assign _T_1116 = _T_1113 != 2'h0;
  assign _T_1117 = _T_1113 | _T_1114;
  assign _T_1118 = _T_1117[1];
  assign _T_1119 = {_T_1116,_T_1118};
  assign _T_1120 = {_T_1111,_T_1119};
  assign _T_1121 = {_T_1106,_T_1120};
  assign _T_1129 = addresses_0_bits == io_r_2_addr;
  assign _T_1130 = addresses_0_valid & _T_1129;
  assign _T_1131 = addresses_1_bits == io_r_2_addr;
  assign _T_1132 = addresses_1_valid & _T_1131;
  assign _T_1133 = addresses_2_bits == io_r_2_addr;
  assign _T_1134 = addresses_2_valid & _T_1133;
  assign _T_1135 = addresses_3_bits == io_r_2_addr;
  assign _T_1136 = addresses_3_valid & _T_1135;
  assign _T_1137 = addresses_4_bits == io_r_2_addr;
  assign _T_1138 = addresses_4_valid & _T_1137;
  assign _T_1139 = addresses_5_bits == io_r_2_addr;
  assign _T_1140 = addresses_5_valid & _T_1139;
  assign _T_1141 = addresses_6_bits == io_r_2_addr;
  assign _T_1142 = addresses_6_valid & _T_1141;
  assign _T_1143 = addresses_7_bits == io_r_2_addr;
  assign _T_1144 = addresses_7_valid & _T_1143;
  assign _T_1145 = addresses_8_bits == io_r_2_addr;
  assign _T_1146 = addresses_8_valid & _T_1145;
  assign _T_1147 = addresses_9_bits == io_r_2_addr;
  assign _T_1148 = addresses_9_valid & _T_1147;
  assign _T_1149 = addresses_10_bits == io_r_2_addr;
  assign _T_1150 = addresses_10_valid & _T_1149;
  assign _T_1151 = addresses_11_bits == io_r_2_addr;
  assign _T_1152 = addresses_11_valid & _T_1151;
  assign _T_1153 = addresses_12_bits == io_r_2_addr;
  assign _T_1154 = addresses_12_valid & _T_1153;
  assign _T_1155 = addresses_13_bits == io_r_2_addr;
  assign _T_1156 = addresses_13_valid & _T_1155;
  assign _T_1157 = addresses_14_bits == io_r_2_addr;
  assign _T_1158 = addresses_14_valid & _T_1157;
  assign _T_1159 = addresses_15_bits == io_r_2_addr;
  assign _T_1160 = addresses_15_valid & _T_1159;
  assign _T_1161 = addresses_16_bits == io_r_2_addr;
  assign _T_1162 = addresses_16_valid & _T_1161;
  assign _T_1163 = addresses_17_bits == io_r_2_addr;
  assign _T_1164 = addresses_17_valid & _T_1163;
  assign _T_1165 = addresses_18_bits == io_r_2_addr;
  assign _T_1166 = addresses_18_valid & _T_1165;
  assign _T_1167 = addresses_19_bits == io_r_2_addr;
  assign _T_1168 = addresses_19_valid & _T_1167;
  assign _T_1169 = addresses_20_bits == io_r_2_addr;
  assign _T_1170 = addresses_20_valid & _T_1169;
  assign _T_1171 = addresses_21_bits == io_r_2_addr;
  assign _T_1172 = addresses_21_valid & _T_1171;
  assign _T_1173 = addresses_22_bits == io_r_2_addr;
  assign _T_1174 = addresses_22_valid & _T_1173;
  assign _T_1175 = addresses_23_bits == io_r_2_addr;
  assign _T_1176 = addresses_23_valid & _T_1175;
  assign _T_1177 = addresses_24_bits == io_r_2_addr;
  assign _T_1178 = addresses_24_valid & _T_1177;
  assign _T_1179 = addresses_25_bits == io_r_2_addr;
  assign _T_1180 = addresses_25_valid & _T_1179;
  assign _T_1181 = addresses_26_bits == io_r_2_addr;
  assign _T_1182 = addresses_26_valid & _T_1181;
  assign _T_1183 = addresses_27_bits == io_r_2_addr;
  assign _T_1184 = addresses_27_valid & _T_1183;
  assign _T_1185 = addresses_28_bits == io_r_2_addr;
  assign _T_1186 = addresses_28_valid & _T_1185;
  assign _T_1187 = addresses_29_bits == io_r_2_addr;
  assign _T_1188 = addresses_29_valid & _T_1187;
  assign _T_1189 = addresses_30_bits == io_r_2_addr;
  assign _T_1190 = addresses_30_valid & _T_1189;
  assign _T_1191 = addresses_31_bits == io_r_2_addr;
  assign _T_1192 = addresses_31_valid & _T_1191;
  assign _T_1230 = {_T_1132,_T_1130};
  assign _T_1231 = {_T_1136,_T_1134};
  assign _T_1232 = {_T_1231,_T_1230};
  assign _T_1233 = {_T_1140,_T_1138};
  assign _T_1234 = {_T_1144,_T_1142};
  assign _T_1235 = {_T_1234,_T_1233};
  assign _T_1236 = {_T_1235,_T_1232};
  assign _T_1237 = {_T_1148,_T_1146};
  assign _T_1238 = {_T_1152,_T_1150};
  assign _T_1239 = {_T_1238,_T_1237};
  assign _T_1240 = {_T_1156,_T_1154};
  assign _T_1241 = {_T_1160,_T_1158};
  assign _T_1242 = {_T_1241,_T_1240};
  assign _T_1243 = {_T_1242,_T_1239};
  assign _T_1244 = {_T_1243,_T_1236};
  assign _T_1245 = {_T_1164,_T_1162};
  assign _T_1246 = {_T_1168,_T_1166};
  assign _T_1247 = {_T_1246,_T_1245};
  assign _T_1248 = {_T_1172,_T_1170};
  assign _T_1249 = {_T_1176,_T_1174};
  assign _T_1250 = {_T_1249,_T_1248};
  assign _T_1251 = {_T_1250,_T_1247};
  assign _T_1252 = {_T_1180,_T_1178};
  assign _T_1253 = {_T_1184,_T_1182};
  assign _T_1254 = {_T_1253,_T_1252};
  assign _T_1255 = {_T_1188,_T_1186};
  assign _T_1256 = {_T_1192,_T_1190};
  assign _T_1257 = {_T_1256,_T_1255};
  assign _T_1258 = {_T_1257,_T_1254};
  assign _T_1259 = {_T_1258,_T_1251};
  assign _T_1260 = {_T_1259,_T_1244};
  assign _T_1262 = _T_1260 != 32'h0;
  assign _T_1263 = _T_1260[31:16];
  assign _T_1264 = _T_1260[15:0];
  assign _T_1266 = _T_1263 != 16'h0;
  assign _T_1267 = _T_1263 | _T_1264;
  assign _T_1268 = _T_1267[15:8];
  assign _T_1269 = _T_1267[7:0];
  assign _T_1271 = _T_1268 != 8'h0;
  assign _T_1272 = _T_1268 | _T_1269;
  assign _T_1273 = _T_1272[7:4];
  assign _T_1274 = _T_1272[3:0];
  assign _T_1276 = _T_1273 != 4'h0;
  assign _T_1277 = _T_1273 | _T_1274;
  assign _T_1278 = _T_1277[3:2];
  assign _T_1279 = _T_1277[1:0];
  assign _T_1281 = _T_1278 != 2'h0;
  assign _T_1282 = _T_1278 | _T_1279;
  assign _T_1283 = _T_1282[1];
  assign _T_1284 = {_T_1281,_T_1283};
  assign _T_1285 = {_T_1276,_T_1284};
  assign _T_1286 = {_T_1271,_T_1285};
  assign _T_1297 = nextAddr + 6'h1;
  assign _T_1298 = _T_1297[5:0];
  assign _T_1463 = _T_932 == 1'h0;
  assign _T_1465 = _T_932 ? {{1'd0}, _GEN_393} : nextAddr;
  assign _GEN_264 = 5'h0 == _GEN_400;
  assign _GEN_265 = 5'h1 == _GEN_400;
  assign _GEN_266 = 5'h2 == _GEN_400;
  assign _GEN_267 = 5'h3 == _GEN_400;
  assign _GEN_268 = 5'h4 == _GEN_400;
  assign _GEN_269 = 5'h5 == _GEN_400;
  assign _GEN_270 = 5'h6 == _GEN_400;
  assign _GEN_271 = 5'h7 == _GEN_400;
  assign _GEN_272 = 5'h8 == _GEN_400;
  assign _GEN_273 = 5'h9 == _GEN_400;
  assign _GEN_274 = 5'ha == _GEN_400;
  assign _GEN_275 = 5'hb == _GEN_400;
  assign _GEN_276 = 5'hc == _GEN_400;
  assign _GEN_277 = 5'hd == _GEN_400;
  assign _GEN_278 = 5'he == _GEN_400;
  assign _GEN_279 = 5'hf == _GEN_400;
  assign _GEN_280 = 5'h10 == _GEN_400;
  assign _GEN_281 = 5'h11 == _GEN_400;
  assign _GEN_282 = 5'h12 == _GEN_400;
  assign _GEN_283 = 5'h13 == _GEN_400;
  assign _GEN_284 = 5'h14 == _GEN_400;
  assign _GEN_285 = 5'h15 == _GEN_400;
  assign _GEN_286 = 5'h16 == _GEN_400;
  assign _GEN_287 = 5'h17 == _GEN_400;
  assign _GEN_288 = 5'h18 == _GEN_400;
  assign _GEN_289 = 5'h19 == _GEN_400;
  assign _GEN_290 = 5'h1a == _GEN_400;
  assign _GEN_291 = 5'h1b == _GEN_400;
  assign _GEN_292 = 5'h1c == _GEN_400;
  assign _GEN_293 = 5'h1d == _GEN_400;
  assign _GEN_294 = 5'h1e == _GEN_400;
  assign _GEN_295 = 5'h1f == _GEN_400;
  assign _T_1488 = _T_1463 ? _T_1298 : nextAddr;
  assign _T_1489 = addresses_0_bits == io_w_1_addr;
  assign _T_1490 = addresses_0_valid & _T_1489;
  assign _T_1491 = addresses_1_bits == io_w_1_addr;
  assign _T_1492 = addresses_1_valid & _T_1491;
  assign _T_1493 = addresses_2_bits == io_w_1_addr;
  assign _T_1494 = addresses_2_valid & _T_1493;
  assign _T_1495 = addresses_3_bits == io_w_1_addr;
  assign _T_1496 = addresses_3_valid & _T_1495;
  assign _T_1497 = addresses_4_bits == io_w_1_addr;
  assign _T_1498 = addresses_4_valid & _T_1497;
  assign _T_1499 = addresses_5_bits == io_w_1_addr;
  assign _T_1500 = addresses_5_valid & _T_1499;
  assign _T_1501 = addresses_6_bits == io_w_1_addr;
  assign _T_1502 = addresses_6_valid & _T_1501;
  assign _T_1503 = addresses_7_bits == io_w_1_addr;
  assign _T_1504 = addresses_7_valid & _T_1503;
  assign _T_1505 = addresses_8_bits == io_w_1_addr;
  assign _T_1506 = addresses_8_valid & _T_1505;
  assign _T_1507 = addresses_9_bits == io_w_1_addr;
  assign _T_1508 = addresses_9_valid & _T_1507;
  assign _T_1509 = addresses_10_bits == io_w_1_addr;
  assign _T_1510 = addresses_10_valid & _T_1509;
  assign _T_1511 = addresses_11_bits == io_w_1_addr;
  assign _T_1512 = addresses_11_valid & _T_1511;
  assign _T_1513 = addresses_12_bits == io_w_1_addr;
  assign _T_1514 = addresses_12_valid & _T_1513;
  assign _T_1515 = addresses_13_bits == io_w_1_addr;
  assign _T_1516 = addresses_13_valid & _T_1515;
  assign _T_1517 = addresses_14_bits == io_w_1_addr;
  assign _T_1518 = addresses_14_valid & _T_1517;
  assign _T_1519 = addresses_15_bits == io_w_1_addr;
  assign _T_1520 = addresses_15_valid & _T_1519;
  assign _T_1521 = addresses_16_bits == io_w_1_addr;
  assign _T_1522 = addresses_16_valid & _T_1521;
  assign _T_1523 = addresses_17_bits == io_w_1_addr;
  assign _T_1524 = addresses_17_valid & _T_1523;
  assign _T_1525 = addresses_18_bits == io_w_1_addr;
  assign _T_1526 = addresses_18_valid & _T_1525;
  assign _T_1527 = addresses_19_bits == io_w_1_addr;
  assign _T_1528 = addresses_19_valid & _T_1527;
  assign _T_1529 = addresses_20_bits == io_w_1_addr;
  assign _T_1530 = addresses_20_valid & _T_1529;
  assign _T_1531 = addresses_21_bits == io_w_1_addr;
  assign _T_1532 = addresses_21_valid & _T_1531;
  assign _T_1533 = addresses_22_bits == io_w_1_addr;
  assign _T_1534 = addresses_22_valid & _T_1533;
  assign _T_1535 = addresses_23_bits == io_w_1_addr;
  assign _T_1536 = addresses_23_valid & _T_1535;
  assign _T_1537 = addresses_24_bits == io_w_1_addr;
  assign _T_1538 = addresses_24_valid & _T_1537;
  assign _T_1539 = addresses_25_bits == io_w_1_addr;
  assign _T_1540 = addresses_25_valid & _T_1539;
  assign _T_1541 = addresses_26_bits == io_w_1_addr;
  assign _T_1542 = addresses_26_valid & _T_1541;
  assign _T_1543 = addresses_27_bits == io_w_1_addr;
  assign _T_1544 = addresses_27_valid & _T_1543;
  assign _T_1545 = addresses_28_bits == io_w_1_addr;
  assign _T_1546 = addresses_28_valid & _T_1545;
  assign _T_1547 = addresses_29_bits == io_w_1_addr;
  assign _T_1548 = addresses_29_valid & _T_1547;
  assign _T_1549 = addresses_30_bits == io_w_1_addr;
  assign _T_1550 = addresses_30_valid & _T_1549;
  assign _T_1551 = addresses_31_bits == io_w_1_addr;
  assign _T_1552 = addresses_31_valid & _T_1551;
  assign _T_1590 = {_T_1492,_T_1490};
  assign _T_1591 = {_T_1496,_T_1494};
  assign _T_1592 = {_T_1591,_T_1590};
  assign _T_1593 = {_T_1500,_T_1498};
  assign _T_1594 = {_T_1504,_T_1502};
  assign _T_1595 = {_T_1594,_T_1593};
  assign _T_1596 = {_T_1595,_T_1592};
  assign _T_1597 = {_T_1508,_T_1506};
  assign _T_1598 = {_T_1512,_T_1510};
  assign _T_1599 = {_T_1598,_T_1597};
  assign _T_1600 = {_T_1516,_T_1514};
  assign _T_1601 = {_T_1520,_T_1518};
  assign _T_1602 = {_T_1601,_T_1600};
  assign _T_1603 = {_T_1602,_T_1599};
  assign _T_1604 = {_T_1603,_T_1596};
  assign _T_1605 = {_T_1524,_T_1522};
  assign _T_1606 = {_T_1528,_T_1526};
  assign _T_1607 = {_T_1606,_T_1605};
  assign _T_1608 = {_T_1532,_T_1530};
  assign _T_1609 = {_T_1536,_T_1534};
  assign _T_1610 = {_T_1609,_T_1608};
  assign _T_1611 = {_T_1610,_T_1607};
  assign _T_1612 = {_T_1540,_T_1538};
  assign _T_1613 = {_T_1544,_T_1542};
  assign _T_1614 = {_T_1613,_T_1612};
  assign _T_1615 = {_T_1548,_T_1546};
  assign _T_1616 = {_T_1552,_T_1550};
  assign _T_1617 = {_T_1616,_T_1615};
  assign _T_1618 = {_T_1617,_T_1614};
  assign _T_1619 = {_T_1618,_T_1611};
  assign _T_1620 = {_T_1619,_T_1604};
  assign _T_1622 = _T_1620 != 32'h0;
  assign _T_1623 = _T_1620[31:16];
  assign _T_1624 = _T_1620[15:0];
  assign _T_1626 = _T_1623 != 16'h0;
  assign _T_1627 = _T_1623 | _T_1624;
  assign _T_1628 = _T_1627[15:8];
  assign _T_1629 = _T_1627[7:0];
  assign _T_1631 = _T_1628 != 8'h0;
  assign _T_1632 = _T_1628 | _T_1629;
  assign _T_1633 = _T_1632[7:4];
  assign _T_1634 = _T_1632[3:0];
  assign _T_1636 = _T_1633 != 4'h0;
  assign _T_1637 = _T_1633 | _T_1634;
  assign _T_1638 = _T_1637[3:2];
  assign _T_1639 = _T_1637[1:0];
  assign _T_1641 = _T_1638 != 2'h0;
  assign _T_1642 = _T_1638 | _T_1639;
  assign _T_1643 = _T_1642[1];
  assign _T_1644 = {_T_1641,_T_1643};
  assign _T_1645 = {_T_1636,_T_1644};
  assign _T_1646 = {_T_1631,_T_1645};
  assign _T_1647 = {_T_1626,_T_1646};
  assign _T_1649 = _T_1622 == 1'h0;
  assign _T_1650 = io_w_1_en & _T_1649;
  assign _T_1651 = _T_1622 ? {{1'd0}, _T_1647} : _T_1488;
  assign _GEN_328 = 5'h0 == _GEN_404;
  assign _GEN_329 = 5'h1 == _GEN_404;
  assign _GEN_330 = 5'h2 == _GEN_404;
  assign _GEN_331 = 5'h3 == _GEN_404;
  assign _GEN_332 = 5'h4 == _GEN_404;
  assign _GEN_333 = 5'h5 == _GEN_404;
  assign _GEN_334 = 5'h6 == _GEN_404;
  assign _GEN_335 = 5'h7 == _GEN_404;
  assign _GEN_336 = 5'h8 == _GEN_404;
  assign _GEN_337 = 5'h9 == _GEN_404;
  assign _GEN_338 = 5'ha == _GEN_404;
  assign _GEN_339 = 5'hb == _GEN_404;
  assign _GEN_340 = 5'hc == _GEN_404;
  assign _GEN_341 = 5'hd == _GEN_404;
  assign _GEN_342 = 5'he == _GEN_404;
  assign _GEN_343 = 5'hf == _GEN_404;
  assign _GEN_344 = 5'h10 == _GEN_404;
  assign _GEN_345 = 5'h11 == _GEN_404;
  assign _GEN_346 = 5'h12 == _GEN_404;
  assign _GEN_347 = 5'h13 == _GEN_404;
  assign _GEN_348 = 5'h14 == _GEN_404;
  assign _GEN_349 = 5'h15 == _GEN_404;
  assign _GEN_350 = 5'h16 == _GEN_404;
  assign _GEN_351 = 5'h17 == _GEN_404;
  assign _GEN_352 = 5'h18 == _GEN_404;
  assign _GEN_353 = 5'h19 == _GEN_404;
  assign _GEN_354 = 5'h1a == _GEN_404;
  assign _GEN_355 = 5'h1b == _GEN_404;
  assign _GEN_356 = 5'h1c == _GEN_404;
  assign _GEN_357 = 5'h1d == _GEN_404;
  assign _GEN_358 = 5'h1e == _GEN_404;
  assign _GEN_359 = 5'h1f == _GEN_404;
  assign _T_1672 = _T_1488 + 6'h1;
  assign _T_1673 = _T_1672[5:0];
  assign nextAddrUpdate = _T_1650 ? _T_1673 : _T_1488;
  assign _T_1675 = nextAddrUpdate <= 6'h20;
  assign _T_1678 = _T_1675 | reset;
  assign _T_1680 = _T_1678 == 1'h0;
  assign io_r_1_data = _T_1097 ? mem__T_1124_data : 32'h0;
  assign io_r_2_data = _T_1262 ? mem__T_1289_data : 32'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  addresses_0_valid = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  addresses_0_bits = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  addresses_1_valid = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  addresses_1_bits = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  addresses_2_valid = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  addresses_2_bits = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  addresses_3_valid = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  addresses_3_bits = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  addresses_4_valid = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  addresses_4_bits = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  addresses_5_valid = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  addresses_5_bits = _RAND_12[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  addresses_6_valid = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  addresses_6_bits = _RAND_14[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  addresses_7_valid = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  addresses_7_bits = _RAND_16[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  addresses_8_valid = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  addresses_8_bits = _RAND_18[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  addresses_9_valid = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  addresses_9_bits = _RAND_20[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  addresses_10_valid = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  addresses_10_bits = _RAND_22[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  addresses_11_valid = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  addresses_11_bits = _RAND_24[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  addresses_12_valid = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  addresses_12_bits = _RAND_26[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  addresses_13_valid = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  addresses_13_bits = _RAND_28[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  addresses_14_valid = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  addresses_14_bits = _RAND_30[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  addresses_15_valid = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  addresses_15_bits = _RAND_32[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  addresses_16_valid = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  addresses_16_bits = _RAND_34[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  addresses_17_valid = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  addresses_17_bits = _RAND_36[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  addresses_18_valid = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  addresses_18_bits = _RAND_38[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  addresses_19_valid = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  addresses_19_bits = _RAND_40[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  addresses_20_valid = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  addresses_20_bits = _RAND_42[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  addresses_21_valid = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  addresses_21_bits = _RAND_44[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  addresses_22_valid = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  addresses_22_bits = _RAND_46[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  addresses_23_valid = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  addresses_23_bits = _RAND_48[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  addresses_24_valid = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  addresses_24_bits = _RAND_50[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  addresses_25_valid = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  addresses_25_bits = _RAND_52[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  addresses_26_valid = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  addresses_26_bits = _RAND_54[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  addresses_27_valid = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  addresses_27_bits = _RAND_56[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  addresses_28_valid = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  addresses_28_bits = _RAND_58[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  addresses_29_valid = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  addresses_29_bits = _RAND_60[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  addresses_30_valid = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  addresses_30_bits = _RAND_62[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  addresses_31_valid = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  addresses_31_bits = _RAND_64[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{$random}};
  nextAddr = _RAND_65[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(mem__T_1484_en & mem__T_1484_mask) begin
      mem[mem__T_1484_addr] <= mem__T_1484_data;
    end
    if(mem__T_1670_en & mem__T_1670_mask) begin
      mem[mem__T_1670_addr] <= mem__T_1670_data;
    end
    if (metaReset) begin
      addresses_0_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_0_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_328) begin
            addresses_0_valid <= 1'h1;
          end else begin
            if (_GEN_264) begin
              addresses_0_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_264) begin
            addresses_0_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_0_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_0_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_328) begin
            addresses_0_bits <= io_w_1_addr;
          end else begin
            if (_GEN_264) begin
              addresses_0_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_264) begin
            addresses_0_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_1_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_1_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_329) begin
            addresses_1_valid <= 1'h1;
          end else begin
            if (_GEN_265) begin
              addresses_1_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_265) begin
            addresses_1_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_1_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_1_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_329) begin
            addresses_1_bits <= io_w_1_addr;
          end else begin
            if (_GEN_265) begin
              addresses_1_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_265) begin
            addresses_1_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_2_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_2_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_330) begin
            addresses_2_valid <= 1'h1;
          end else begin
            if (_GEN_266) begin
              addresses_2_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_266) begin
            addresses_2_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_2_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_2_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_330) begin
            addresses_2_bits <= io_w_1_addr;
          end else begin
            if (_GEN_266) begin
              addresses_2_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_266) begin
            addresses_2_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_3_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_3_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_331) begin
            addresses_3_valid <= 1'h1;
          end else begin
            if (_GEN_267) begin
              addresses_3_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_267) begin
            addresses_3_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_3_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_3_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_331) begin
            addresses_3_bits <= io_w_1_addr;
          end else begin
            if (_GEN_267) begin
              addresses_3_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_267) begin
            addresses_3_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_4_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_4_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_332) begin
            addresses_4_valid <= 1'h1;
          end else begin
            if (_GEN_268) begin
              addresses_4_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_268) begin
            addresses_4_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_4_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_4_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_332) begin
            addresses_4_bits <= io_w_1_addr;
          end else begin
            if (_GEN_268) begin
              addresses_4_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_268) begin
            addresses_4_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_5_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_5_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_333) begin
            addresses_5_valid <= 1'h1;
          end else begin
            if (_GEN_269) begin
              addresses_5_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_269) begin
            addresses_5_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_5_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_5_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_333) begin
            addresses_5_bits <= io_w_1_addr;
          end else begin
            if (_GEN_269) begin
              addresses_5_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_269) begin
            addresses_5_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_6_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_6_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_334) begin
            addresses_6_valid <= 1'h1;
          end else begin
            if (_GEN_270) begin
              addresses_6_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_270) begin
            addresses_6_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_6_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_6_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_334) begin
            addresses_6_bits <= io_w_1_addr;
          end else begin
            if (_GEN_270) begin
              addresses_6_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_270) begin
            addresses_6_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_7_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_7_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_335) begin
            addresses_7_valid <= 1'h1;
          end else begin
            if (_GEN_271) begin
              addresses_7_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_271) begin
            addresses_7_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_7_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_7_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_335) begin
            addresses_7_bits <= io_w_1_addr;
          end else begin
            if (_GEN_271) begin
              addresses_7_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_271) begin
            addresses_7_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_8_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_8_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_336) begin
            addresses_8_valid <= 1'h1;
          end else begin
            if (_GEN_272) begin
              addresses_8_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_272) begin
            addresses_8_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_8_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_8_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_336) begin
            addresses_8_bits <= io_w_1_addr;
          end else begin
            if (_GEN_272) begin
              addresses_8_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_272) begin
            addresses_8_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_9_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_9_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_337) begin
            addresses_9_valid <= 1'h1;
          end else begin
            if (_GEN_273) begin
              addresses_9_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_273) begin
            addresses_9_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_9_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_9_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_337) begin
            addresses_9_bits <= io_w_1_addr;
          end else begin
            if (_GEN_273) begin
              addresses_9_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_273) begin
            addresses_9_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_10_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_10_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_338) begin
            addresses_10_valid <= 1'h1;
          end else begin
            if (_GEN_274) begin
              addresses_10_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_274) begin
            addresses_10_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_10_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_10_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_338) begin
            addresses_10_bits <= io_w_1_addr;
          end else begin
            if (_GEN_274) begin
              addresses_10_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_274) begin
            addresses_10_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_11_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_11_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_339) begin
            addresses_11_valid <= 1'h1;
          end else begin
            if (_GEN_275) begin
              addresses_11_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_275) begin
            addresses_11_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_11_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_11_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_339) begin
            addresses_11_bits <= io_w_1_addr;
          end else begin
            if (_GEN_275) begin
              addresses_11_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_275) begin
            addresses_11_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_12_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_12_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_340) begin
            addresses_12_valid <= 1'h1;
          end else begin
            if (_GEN_276) begin
              addresses_12_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_276) begin
            addresses_12_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_12_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_12_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_340) begin
            addresses_12_bits <= io_w_1_addr;
          end else begin
            if (_GEN_276) begin
              addresses_12_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_276) begin
            addresses_12_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_13_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_13_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_341) begin
            addresses_13_valid <= 1'h1;
          end else begin
            if (_GEN_277) begin
              addresses_13_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_277) begin
            addresses_13_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_13_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_13_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_341) begin
            addresses_13_bits <= io_w_1_addr;
          end else begin
            if (_GEN_277) begin
              addresses_13_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_277) begin
            addresses_13_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_14_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_14_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_342) begin
            addresses_14_valid <= 1'h1;
          end else begin
            if (_GEN_278) begin
              addresses_14_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_278) begin
            addresses_14_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_14_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_14_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_342) begin
            addresses_14_bits <= io_w_1_addr;
          end else begin
            if (_GEN_278) begin
              addresses_14_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_278) begin
            addresses_14_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_15_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_15_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_343) begin
            addresses_15_valid <= 1'h1;
          end else begin
            if (_GEN_279) begin
              addresses_15_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_279) begin
            addresses_15_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_15_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_15_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_343) begin
            addresses_15_bits <= io_w_1_addr;
          end else begin
            if (_GEN_279) begin
              addresses_15_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_279) begin
            addresses_15_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_16_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_16_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_344) begin
            addresses_16_valid <= 1'h1;
          end else begin
            if (_GEN_280) begin
              addresses_16_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_280) begin
            addresses_16_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_16_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_16_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_344) begin
            addresses_16_bits <= io_w_1_addr;
          end else begin
            if (_GEN_280) begin
              addresses_16_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_280) begin
            addresses_16_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_17_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_17_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_345) begin
            addresses_17_valid <= 1'h1;
          end else begin
            if (_GEN_281) begin
              addresses_17_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_281) begin
            addresses_17_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_17_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_17_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_345) begin
            addresses_17_bits <= io_w_1_addr;
          end else begin
            if (_GEN_281) begin
              addresses_17_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_281) begin
            addresses_17_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_18_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_18_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_346) begin
            addresses_18_valid <= 1'h1;
          end else begin
            if (_GEN_282) begin
              addresses_18_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_282) begin
            addresses_18_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_18_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_18_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_346) begin
            addresses_18_bits <= io_w_1_addr;
          end else begin
            if (_GEN_282) begin
              addresses_18_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_282) begin
            addresses_18_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_19_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_19_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_347) begin
            addresses_19_valid <= 1'h1;
          end else begin
            if (_GEN_283) begin
              addresses_19_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_283) begin
            addresses_19_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_19_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_19_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_347) begin
            addresses_19_bits <= io_w_1_addr;
          end else begin
            if (_GEN_283) begin
              addresses_19_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_283) begin
            addresses_19_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_20_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_20_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_348) begin
            addresses_20_valid <= 1'h1;
          end else begin
            if (_GEN_284) begin
              addresses_20_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_284) begin
            addresses_20_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_20_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_20_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_348) begin
            addresses_20_bits <= io_w_1_addr;
          end else begin
            if (_GEN_284) begin
              addresses_20_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_284) begin
            addresses_20_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_21_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_21_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_349) begin
            addresses_21_valid <= 1'h1;
          end else begin
            if (_GEN_285) begin
              addresses_21_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_285) begin
            addresses_21_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_21_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_21_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_349) begin
            addresses_21_bits <= io_w_1_addr;
          end else begin
            if (_GEN_285) begin
              addresses_21_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_285) begin
            addresses_21_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_22_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_22_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_350) begin
            addresses_22_valid <= 1'h1;
          end else begin
            if (_GEN_286) begin
              addresses_22_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_286) begin
            addresses_22_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_22_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_22_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_350) begin
            addresses_22_bits <= io_w_1_addr;
          end else begin
            if (_GEN_286) begin
              addresses_22_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_286) begin
            addresses_22_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_23_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_23_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_351) begin
            addresses_23_valid <= 1'h1;
          end else begin
            if (_GEN_287) begin
              addresses_23_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_287) begin
            addresses_23_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_23_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_23_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_351) begin
            addresses_23_bits <= io_w_1_addr;
          end else begin
            if (_GEN_287) begin
              addresses_23_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_287) begin
            addresses_23_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_24_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_24_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_352) begin
            addresses_24_valid <= 1'h1;
          end else begin
            if (_GEN_288) begin
              addresses_24_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_288) begin
            addresses_24_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_24_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_24_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_352) begin
            addresses_24_bits <= io_w_1_addr;
          end else begin
            if (_GEN_288) begin
              addresses_24_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_288) begin
            addresses_24_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_25_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_25_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_353) begin
            addresses_25_valid <= 1'h1;
          end else begin
            if (_GEN_289) begin
              addresses_25_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_289) begin
            addresses_25_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_25_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_25_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_353) begin
            addresses_25_bits <= io_w_1_addr;
          end else begin
            if (_GEN_289) begin
              addresses_25_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_289) begin
            addresses_25_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_26_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_26_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_354) begin
            addresses_26_valid <= 1'h1;
          end else begin
            if (_GEN_290) begin
              addresses_26_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_290) begin
            addresses_26_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_26_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_26_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_354) begin
            addresses_26_bits <= io_w_1_addr;
          end else begin
            if (_GEN_290) begin
              addresses_26_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_290) begin
            addresses_26_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_27_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_27_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_355) begin
            addresses_27_valid <= 1'h1;
          end else begin
            if (_GEN_291) begin
              addresses_27_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_291) begin
            addresses_27_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_27_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_27_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_355) begin
            addresses_27_bits <= io_w_1_addr;
          end else begin
            if (_GEN_291) begin
              addresses_27_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_291) begin
            addresses_27_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_28_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_28_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_356) begin
            addresses_28_valid <= 1'h1;
          end else begin
            if (_GEN_292) begin
              addresses_28_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_292) begin
            addresses_28_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_28_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_28_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_356) begin
            addresses_28_bits <= io_w_1_addr;
          end else begin
            if (_GEN_292) begin
              addresses_28_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_292) begin
            addresses_28_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_29_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_29_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_357) begin
            addresses_29_valid <= 1'h1;
          end else begin
            if (_GEN_293) begin
              addresses_29_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_293) begin
            addresses_29_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_29_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_29_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_357) begin
            addresses_29_bits <= io_w_1_addr;
          end else begin
            if (_GEN_293) begin
              addresses_29_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_293) begin
            addresses_29_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_30_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_30_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_358) begin
            addresses_30_valid <= 1'h1;
          end else begin
            if (_GEN_294) begin
              addresses_30_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_294) begin
            addresses_30_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_30_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_30_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_358) begin
            addresses_30_bits <= io_w_1_addr;
          end else begin
            if (_GEN_294) begin
              addresses_30_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_294) begin
            addresses_30_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_31_valid <= 1'h0;
    end else begin
      if (reset) begin
        addresses_31_valid <= 1'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_359) begin
            addresses_31_valid <= 1'h1;
          end else begin
            if (_GEN_295) begin
              addresses_31_valid <= 1'h1;
            end
          end
        end else begin
          if (_GEN_295) begin
            addresses_31_valid <= 1'h1;
          end
        end
      end
    end
    if (metaReset) begin
      addresses_31_bits <= 5'h0;
    end else begin
      if (reset) begin
        addresses_31_bits <= 5'h0;
      end else begin
        if (io_w_1_en) begin
          if (_GEN_359) begin
            addresses_31_bits <= io_w_1_addr;
          end else begin
            if (_GEN_295) begin
              addresses_31_bits <= 5'h0;
            end
          end
        end else begin
          if (_GEN_295) begin
            addresses_31_bits <= 5'h0;
          end
        end
      end
    end
    if (metaReset) begin
      nextAddr <= 6'h0;
    end else begin
      if (reset) begin
        nextAddr <= 6'h0;
      end else begin
        if (_T_1650) begin
          nextAddr <= _T_1673;
        end else begin
          if (_T_1463) begin
            nextAddr <= _T_1298;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1680) begin
          $fwrite(32'h80000002,"Assertion failed: SparseMem ran out of space with size %d, increase size in ReplaceMemsTransform!\n    at SparseMem.scala:103 assert(nextAddrUpdate <= depth.U,\n",6'h20);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1680) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Core( // @[:Sodor3Stage.fir@3688.2]
  input         metaReset,
  input         clock, // @[:Sodor3Stage.fir@3689.4]
  input         reset, // @[:Sodor3Stage.fir@3690.4]
  output [31:0] io_imem_req_bits_addr, // @[:Sodor3Stage.fir@3691.4]
  input  [31:0] io_imem_resp_bits_data, // @[:Sodor3Stage.fir@3691.4]
  output [31:0] io_dmem_req_bits_addr, // @[:Sodor3Stage.fir@3691.4]
  output [31:0] io_dmem_req_bits_data, // @[:Sodor3Stage.fir@3691.4]
  output        io_dmem_req_bits_fcn, // @[:Sodor3Stage.fir@3691.4]
  output [2:0]  io_dmem_req_bits_typ, // @[:Sodor3Stage.fir@3691.4]
  input  [31:0] io_dmem_resp_bits_data, // @[:Sodor3Stage.fir@3691.4]
  output        _GEN_338,
  output        _GEN_224,
  output        _GEN_218,
  output        _GEN_21,
  output        _GEN_91,
  output        _GEN_323,
  output        _GEN_302,
  output        _GEN_51,
  output        _GEN_304,
  output        _GEN_199,
  output        _GEN_6,
  output        _GEN_148,
  output        _GEN_239,
  output        _GEN_403,
  output        _GEN_1,
  output        _GEN_24,
  output        _GEN_247,
  output        _GEN_106,
  output        _GEN_317,
  output        _GEN_133,
  output        _GEN_205,
  output        _GEN_385,
  output        _GEN_39,
  output        _GEN_232,
  output        _GEN_418,
  output        _GEN_127,
  output        _GEN_197,
  output        _GEN_331,
  output        _GEN_190,
  output        _GEN_12,
  output        _GEN_226,
  output        _GEN_296,
  output        _GEN_9_0,
  output        _GEN_45,
  output        _GEN_112,
  output        _GEN_298,
  output        _GEN_203,
  output        _GEN_72,
  output        _GEN_211,
  output        _GEN_325,
  output        _GEN_397,
  output        _GEN_0,
  output        _GEN_424,
  output        _GEN_30,
  output        _GEN_310,
  output        _GEN_319,
  output        _GEN_66,
  output        _GEN_9_1,
  output        _GEN_212,
  output        _GEN_220,
  output        _GEN_214,
  output        _GEN_100,
  output        _GEN_109,
  output        _GEN_320,
  output        _GEN_313,
  output        _GEN_282,
  output        _GEN_200,
  output        _GEN_177,
  output        _GEN_208,
  output        _GEN_388,
  output        _GEN_391,
  output        _GEN_381,
  output        _GEN_412,
  output        _GEN_27,
  output        _GEN_276,
  output        _GEN_191,
  output        _GEN_181,
  output        _GEN_54,
  output        _GEN_193,
  output        _GEN_190_0,
  output        _GEN_15,
  output        _GEN_289,
  output        _GEN_12_0,
  output        _GEN_406,
  output        _GEN_299,
  output        _GEN_48,
  output        _GEN_115,
  output        _GEN_311,
  output        _GEN_206,
  output        _GEN_367,
  output        _GEN_175,
  output        _GEN_6_0,
  output        _GEN_305,
  output        _GEN_33,
  output        _GEN_274,
  output        _GEN_121,
  output        _GEN_307,
  output        _GEN_373,
  output        _GEN_375,
  output        _GEN_229,
  output        _GEN_94,
  output        _GEN_292,
  output        _GEN_183,
  output        _GEN_376,
  output        _GEN_382,
  output        _GEN_0_0,
  output        _GEN_10,
  output        _GEN_370,
  output        _GEN_349,
  output        _GEN_196,
  output        _GEN_186,
  output        _GEN_262,
  output        _GEN_400,
  output        _GEN_103,
  output        _GEN_264,
  output        _GEN_295,
  output        _GEN_355,
  output        _GEN_159,
  output        _GEN_202,
  output        _GEN_171,
  output        _GEN_357,
  output        _GEN_270,
  output        _GEN_277,
  output        _GEN_384,
  output        _GEN_36,
  output        _GEN_285,
  output        _GEN_165,
  output        _GEN_279,
  output        _GEN_194,
  output        _GEN_184,
  output        _GEN_378,
  output        _GEN_293,
  output        _GEN_21_0,
  output        _GEN_301,
  output        _GEN_157,
  output        _GEN_3_0,
  output        _GEN_361,
  output        _GEN_394,
  output        _GEN_15_0,
  output        _GEN_256,
  output        _GEN_363,
  output        _GEN_9_2,
  output        _GEN_258,
  output        _GEN_97,
  output        _GEN_283,
  output        _GEN_163,
  output        _GEN_178,
  output        _GEN_345,
  output        _GEN_339,
  output        _GEN_8,
  output        _GEN_11,
  output        _GEN_18,
  output        _GEN_259,
  output        _GEN_147,
  output        _GEN_358,
  output        _GEN_330,
  output        _GEN_172,
  output        _GEN_86,
  output        _GEN_13,
  output        _GEN_271,
  output        _GEN_265,
  output        _GEN_280,
  output        _GEN_160,
  output        _GEN_273,
  output        _GEN_343,
  output        _GEN_379,
  output        _GEN_351,
  output        _GEN_238,
  output        _GEN_231,
  output        _GEN_189,
  output        _GEN_337,
  output        _GEN_153,
  output        _GEN_288,
  output        _GEN_364,
  output        _GEN_244,
  output        _GEN_366,
  output        _GEN_252,
  output        _GEN_180,
  output        _GEN_166,
  output        _GEN_71,
  output        _GEN_174,
  output        _GEN_168,
  output        _GEN_372,
  output        _GEN_3_1,
  output        _GEN_387,
  output        _GEN_246,
  output        _GEN_267,
  output        _GEN_286,
  output        _GEN_151,
  output        _GEN_187,
  output        _GEN_354,
  output        _GEN_213,
  output        _GEN_249,
  output        _GEN_319_0,
  output        _GEN_268,
  output        _GEN_240,
  output        _GEN_141,
  output        _GEN_135,
  output        _GEN_226_0,
  output        _GEN_234,
  output        _GEN_348,
  output        _GEN_261,
  output        _GEN_312,
  output        _GEN_53,
  output        _GEN_333,
  output        _GEN_147_0,
  output        _GEN_68,
  output        _GEN_156,
  output        _GEN_352,
  output        _GEN_247_0,
  output        _GEN_360,
  output        _GEN_369,
  output        _GEN_325_0,
  output        _GEN_2,
  output        _GEN_74,
  output        _GEN_327,
  output        _GEN_169,
  output        _GEN_89,
  output        _GEN_162,
  output        _GEN_232_0,
  output        _GEN_426,
  output        _GEN_7_0,
  output        _GEN_331_0,
  output        _GEN_129,
  output        _GEN_346,
  output        _GEN_154,
  output        _GEN_340,
  output        _GEN_253,
  output        _GEN_228,
  output        _GEN_411,
  output        _GEN_255,
  output        _GEN_120,
  output        _GEN_211_0,
  output        _GEN_80,
  output        _GEN_220_0,
  output        _GEN_342,
  output        _GEN_229_0,
  output        _GEN_393,
  output        _GEN_292_0,
  output        _GEN_307_0,
  output        _GEN_193_0,
  output        _GEN_56,
  output        _GEN_144,
  output        _GEN_17,
  output        _GEN_11_1,
  output        _GEN_408,
  output        _GEN_222,
  output        _GEN_313_0,
  output        _GEN_117,
  output        _GEN_328,
  output        _GEN_321,
  output        _GEN_2_0,
  output        _GEN_235,
  output        _GEN_243,
  output        _GEN_237,
  output        _GEN_123,
  output        _GEN_102,
  output        _GEN_3_2,
  output        _GEN_62,
  output        _GEN_150,
  output        _GEN_336,
  output        _GEN_201,
  output        _GEN_195,
  output        _GEN_23,
  output        _GEN_414,
  output        _GEN_250,
  output        _GEN_300,
  output        _GEN_294,
  output        _GEN_309,
  output        _GEN_77,
  output        _GEN_208_0,
  output        _GEN_83,
  output        _GEN_214_0,
  output        _GEN_216,
  output        _GEN_241,
  output        _GEN_420,
  output        _GEN_35,
  output        _GEN_5_0,
  output        _GEN_41,
  output        _GEN_315,
  output        _GEN_429,
  output        _GEN_138,
  output        _GEN_334,
  output        _GEN_217,
  output        _GEN_402,
  output        _GEN_17_0,
  output        _GEN_225,
  output        _GEN_105,
  output        _GEN_316,
  output        _GEN_50,
  output        _GEN_44,
  output        _GEN_324,
  output        _GEN_180_0,
  output        _GEN_318,
  output        _GEN_384_0,
  output        _GEN_396,
  output        _GEN_386,
  output        _GEN_38,
  output        _GEN_301_0,
  output        _GEN_196_0,
  output        _GEN_186_0,
  output        _GEN_65,
  output        _GEN_295_0,
  output        _GEN_20,
  output        _GEN_223,
  output        _GEN_23_0,
  output        _GEN_417,
  output        _GEN_111,
  output        _GEN_322,
  output        _GEN_210,
  output        _GEN_5_1,
  output        _GEN_219,
  output        _GEN_279_0,
  output        _GEN_310_0,
  output        _GEN_285_0,
  output        _GEN_423,
  output        _GEN_132,
  output        _GEN_126,
  output        _GEN_287,
  output        _GEN_202_0,
  output        _GEN_378_0,
  output        _GEN_90,
  output        _GEN_204,
  output        _GEN_99,
  output        _GEN_303,
  output        _GEN_297,
  output        _GEN_59,
  output        _GEN_188,
  output        _GEN_198,
  output        _GEN_351_0,
  output        _GEN_176,
  output        _GEN_387_0,
  output        _GEN_11_2,
  output        _GEN_380,
  output        _GEN_93,
  output        _GEN_161,
  output        _GEN_192,
  output        _GEN_189_0,
  output        _GEN_14_0,
  output        _GEN_372_0,
  output        _GEN_207,
  output        _GEN_267_0,
  output        _GEN_405,
  output        _GEN_260,
  output        _GEN_26,
  output        _GEN_114,
  output        _GEN_269,
  output        _GEN_174_0,
  output        _GEN_205_0,
  output        _GEN_182,
  output        _GEN_399,
  output        _GEN_368,
  output        _GEN_273_0,
  output        _GEN_390,
  output        _GEN_32,
  output        _GEN_281,
  output        _GEN_275,
  output        _GEN_291,
  output        _GEN_168_0,
  output        _GEN_47,
  output        _GEN_199_0,
  output        _GEN_5_2,
  output        _GEN_389,
  output        _GEN_298_0,
  output        _GEN_304_0,
  output        _GEN_306,
  output        _GEN_366_0,
  output        _GEN_8_1,
  output        _GEN_374,
  output        _GEN_108,
  output        _GEN_360_0,
  output        _GEN_288_0,
  output        _GEN_356,
  output        _GEN_375_0,
  output        _GEN_255_0,
  output        _GEN_261_0,
  output        _GEN_20_0,
  output        _GEN_14_1,
  output        _GEN_29,
  output        _GEN_270_0,
  output        _GEN_150_0,
  output        _GEN_333_0,
  output        _GEN_82,
  output        _GEN_177_0,
  output        _GEN_170,
  output        _GEN_381_0,
  output        _GEN_185,
  output        _GEN_1_1,
  output        _GEN_276_0,
  output        _GEN_10_0,
  output        _GEN_278,
  output        _GEN_143,
  output        _GEN_354_0,
  output        _GEN_348_0,
  output        _GEN_249_0,
  output        _GEN_96,
  output        _GEN_9_3,
  output        _GEN_263,
  output        _GEN_164,
  output        _GEN_158,
  output        _GEN_369_0,
  output        _GEN_183_0,
  output        _GEN_362,
  output        _GEN_377,
  output        _GEN_257,
  output        _GEN_282_0,
  output        _GEN_284,
  output        _GEN_179,
  output        _GEN_383,
  output        _GEN_242,
  output        _GEN_8_2,
  output        _GEN_162_0,
  output        _GEN_156_0,
  output        _GEN_341,
  output        _GEN_76,
  output        _GEN_165_0,
  output        _GEN_173,
  output        _GEN_224_0,
  output        _GEN_359,
  output        _GEN_251,
  output        _GEN_131,
  output        _GEN_7_1,
  output        _GEN_146,
  output        _GEN_342_0,
  output        _GEN_350,
  output        _GEN_344,
  output        _GEN_239_0,
  output        _GEN_264_0,
  output        _GEN_272,
  output        _GEN_64,
  output        _GEN_58,
  output        _GEN_159_0,
  output        _GEN_222_0,
  output        _GEN_363_0,
  output        _GEN_357_0,
  output        _GEN_230,
  output        _GEN_365,
  output        _GEN_321_0,
  output        _GEN_7_2,
  output        _GEN_330_0,
  output        _GEN_323_0,
  output        _GEN_85,
  output        _GEN_338_0,
  output        _GEN_79,
  output        _GEN_243_0,
  output        _GEN_2_2,
  output        _GEN_237_0,
  output        _GEN_245,
  output        _GEN_12_1,
  output        _GEN_315_0,
  output        _GEN_336_0,
  output        _GEN_70,
  output        _GEN_152,
  output        _GEN_167,
  output        _GEN_422,
  output        _GEN_258_0,
  output        _GEN_371,
  output        _GEN_266,
  output        _GEN_125,
  output        _GEN_171_0,
  output        _GEN_212_0,
  output        _GEN_303_0,
  output        _GEN_254,
  output        _GEN_146_0,
  output        _GEN_13_0,
  output        _GEN_155,
  output        _GEN_149,
  output        _GEN_225_0,
  output        _GEN_227,
  output        _GEN_113,
  output        _GEN_140,
  output        _GEN_326,
  output        _GEN_7_3,
  output        _GEN_231_0,
  output        _GEN_425,
  output        _GEN_404,
  output        _GEN_240_0,
  output        _GEN_353,
  output        _GEN_248,
  output        _GEN_107,
  output        _GEN_6_3,
  output        _GEN_311_0,
  output        _GEN_339_0,
  output        _GEN_153_0,
  output        _GEN_73,
  output        _GEN_67,
  output        _GEN_347,
  output        _GEN_206_0,
  output        _GEN_252_0,
  output        _GEN_410,
  output        _GEN_297_0,
  output        _GEN_419,
  output        _GEN_233,
  output        _GEN_305_0,
  output        _GEN_128,
  output        _GEN_324_0,
  output        _GEN_332,
  output        _GEN_219_0,
  output        _GEN_88,
  output        _GEN_1_3,
  output        _GEN_246_0,
  output        _GEN_318_0,
  output        _GEN_52,
  output        _GEN_46,
  output        _GEN_134,
  output        _GEN_345_0,
  output        _GEN_204_0,
  output        _GEN_213_0,
  output        _GEN_228_0,
  output        _GEN_221,
  output        _GEN_407,
  output        _GEN_382_0,
  output        _GEN_28,
  output        _GEN_281_0,
  output        _GEN_4_1,
  output        _GEN_40,
  output        _GEN_55,
  output        _GEN_329,
  output        _GEN_194_0,
  output        _GEN_392,
  output        _GEN_0_2,
  output        _GEN_234_0,
  output        _GEN_10_2,
  output        _GEN_236,
  output        _GEN_101,
  output        _GEN_312_0,
  output        _GEN_192_0,
  output        _GEN_306_0,
  output        _GEN_61,
  output        _GEN_207_0,
  output        _GEN_16,
  output        _GEN_22,
  output        _GEN_300_0,
  output        _GEN_34,
  output        _GEN_116,
  output        _GEN_122,
  output        _GEN_327_0,
  output        _GEN_182_0,
  output        _GEN_320_0,
  output        _GEN_215,
  output        _GEN_335,
  output        _GEN_291_0,
  output        _GEN_290,
  output        _GEN_293_0,
  output        _GEN_428,
  output        _GEN_49,
  output        _GEN_137,
  output        _GEN_200_0,
  output        _GEN_209,
  output        _GEN_95,
  output        _GEN_413,
  output        _GEN_314,
  output        _GEN_308,
  output        _GEN_4_2,
  output        _GEN_383_0,
  output        _GEN_16_0,
  output        _GEN_395,
  output        _GEN_385_0,
  output        _GEN_104,
  output        _GEN_195_0,
  output        _GEN_302_0,
  output        _GEN_317_0,
  output        _GEN_203_0,
  output        _GEN_172_0,
  output        _GEN_197_0,
  output        _GEN_370_0,
  output        _GEN_416,
  output        _GEN_22_0,
  output        _GEN_271_0,
  output        _GEN_119,
  output        _GEN_185_0,
  output        _GEN_179_0,
  output        _GEN_216_0,
  output        _GEN_379_0,
  output        _GEN_187_0,
  output        _GEN_401,
  output        _GEN_43,
  output        _GEN_278_0,
  output        _GEN_296_0,
  output        _GEN_286_0,
  output        _GEN_201_0,
  output        _GEN_364_0,
  output        _GEN_1_4,
  output        _GEN_210_0,
  output        _GEN_98,
  output        _GEN_263_0,
  output        _GEN_309_0,
  output        _GEN_37,
  output        _GEN_164_0,
  output        _GEN_110,
  output        _GEN_362_0,
  output        _GEN_19,
  output        _GEN_377_0,
  output        _GEN_218_0,
  output        _GEN_294_0,
  output        _GEN_284_0,
  output        _GEN_371_0,
  output        _GEN_260_0,
  output        _GEN_266_0,
  output        _GEN_380_0,
  output        _GEN_25,
  output        _GEN_365_0,
  output        _GEN_181_0,
  output        _GEN_175_0,
  output        _GEN_251_0,
  output        _GEN_15_1,
  output        _GEN_289_0,
  output        _GEN_359_0,
  output        _GEN_352_0,
  output        _GEN_14_2,
  output        _GEN_152_0,
  output        _GEN_31,
  output        _GEN_274_0,
  output        _GEN_160_0,
  output        _GEN_169_0,
  output        _GEN_191_0,
  output        _GEN_188_0,
  output        _GEN_373_0,
  output        _GEN_19_0,
  output        _GEN_367_0,
  output        _GEN_268_0,
  output        _GEN_173_0,
  output        _GEN_290_0,
  output        _GEN_280_0,
  output        _GEN_287_0,
  output        _GEN_154_0,
  output        _GEN_87,
  output        _GEN_299_0,
  output        _GEN_386_0,
  output        _GEN_10_3,
  output        _GEN_245_0,
  output        _GEN_398,
  output        _GEN_4_3,
  output        _GEN_388_0,
  output        _GEN_253_0,
  output        _GEN_92,
  output        _GEN_5_3,
  output        _GEN_272_0,
  output        _GEN_344_0,
  output        _GEN_198_0,
  output        _GEN_167_0,
  output        _GEN_346_0,
  output        _GEN_334_0,
  output        _GEN_340_0,
  output        _GEN_254_0,
  output        _GEN_13_2,
  output        _GEN_3_4,
  output        _GEN_256_0,
  output        _GEN_328_0,
  output        _GEN_161_0,
  output        _GEN_347_0,
  output        _GEN_81,
  output        _GEN_355_0,
  output        _GEN_170_0,
  output        _GEN_7_5,
  output        _GEN_8_3,
  output        _GEN_275_0,
  output        _GEN_269_0,
  output        _GEN_155_0,
  output        _GEN_277_0,
  output        _GEN_69,
  output        _GEN_157_0,
  output        _GEN_368_0,
  output        _GEN_233_0,
  output        _GEN_227_0,
  output        _GEN_235_0,
  output        _GEN_184_0,
  output        _GEN_326_0,
  output        _GEN_149_0,
  output        _GEN_60,
  output        _GEN_283_0,
  output        _GEN_142,
  output        _GEN_353_0,
  output        _GEN_178_0,
  output        _GEN_248_0,
  output        _GEN_241_0,
  output        _GEN_361_0,
  output        _GEN_136,
  output        _GEN_75,
  output        _GEN_163_0,
  output        _GEN_349_0,
  output        _GEN_374_0,
  output        _GEN_427,
  output        _GEN_376_0,
  output        _GEN_262_0,
  output        _GEN_332_0,
  output        _GEN_176_0,
  output        _GEN_166_0,
  output        _GEN_358_0,
  output        _GEN_314_0,
  output        _GEN_308_0,
  output        _GEN_42,
  output        _GEN_265_0,
  output        _GEN_316_0,
  output        _GEN_130,
  output        _GEN_124,
  output        _GEN_341_0,
  output        _GEN_343_0,
  output        _GEN_223_0,
  output        _GEN_238_0,
  output        _GEN_118,
  output        _GEN_5_4,
  output        _GEN_151_0,
  output        _GEN_145,
  output        _GEN_337_0,
  output        _GEN_18_0,
  output        _GEN_356_0,
  output        _GEN_244_0,
  output        _GEN_409,
  output        _GEN_11_3,
  output        _GEN_322_0,
  output        _GEN_158_0,
  output        _GEN_209_0,
  output        _GEN_78,
  output        _GEN_217_0,
  output        _GEN_221_0,
  output        _GEN_236_0,
  output        _GEN_421,
  output        _GEN_415,
  output        _GEN_335_0,
  output        _GEN_329_0,
  output        _GEN_63,
  output        _GEN_230_0,
  output        _GEN_242_0,
  output        _GEN_257_0,
  output        _GEN_6_4,
  output        _GEN_57,
  output        _GEN_250_0,
  output        _GEN_259_0,
  output        _GEN_139,
  output        _GEN_350_0,
  output        _GEN_215_0,
  output        _GEN_84
);
  wire  frontend_metaReset; // @[core.scala 25:25:Sodor3Stage.fir@3693.4]
  wire  frontend_clock; // @[core.scala 25:25:Sodor3Stage.fir@3693.4]
  wire  frontend_reset; // @[core.scala 25:25:Sodor3Stage.fir@3693.4]
  wire  frontend_io_cpu_req_valid; // @[core.scala 25:25:Sodor3Stage.fir@3693.4]
  wire [31:0] frontend_io_cpu_req_bits_pc; // @[core.scala 25:25:Sodor3Stage.fir@3693.4]
  wire  frontend_io_cpu_resp_ready; // @[core.scala 25:25:Sodor3Stage.fir@3693.4]
  wire  frontend_io_cpu_resp_valid; // @[core.scala 25:25:Sodor3Stage.fir@3693.4]
  wire [31:0] frontend_io_cpu_resp_bits_pc; // @[core.scala 25:25:Sodor3Stage.fir@3693.4]
  wire [31:0] frontend_io_cpu_resp_bits_inst; // @[core.scala 25:25:Sodor3Stage.fir@3693.4]
  wire [31:0] frontend_io_imem_req_bits_addr; // @[core.scala 25:25:Sodor3Stage.fir@3693.4]
  wire [31:0] frontend_io_imem_resp_bits_data; // @[core.scala 25:25:Sodor3Stage.fir@3693.4]
  wire  frontend__GEN_1_0; // @[core.scala 25:25:Sodor3Stage.fir@3693.4]
  wire  frontend__GEN_10_0; // @[core.scala 25:25:Sodor3Stage.fir@3693.4]
  wire  frontend__GEN_13_0; // @[core.scala 25:25:Sodor3Stage.fir@3693.4]
  wire  frontend__GEN_7_1; // @[core.scala 25:25:Sodor3Stage.fir@3693.4]
  wire  frontend__GEN_9_4; // @[core.scala 25:25:Sodor3Stage.fir@3693.4]
  wire  frontend__GEN_12_2; // @[core.scala 25:25:Sodor3Stage.fir@3693.4]
  wire  frontend__GEN_6_4; // @[core.scala 25:25:Sodor3Stage.fir@3693.4]
  wire  frontend__GEN_14_3; // @[core.scala 25:25:Sodor3Stage.fir@3693.4]
  wire  frontend__GEN_5_4; // @[core.scala 25:25:Sodor3Stage.fir@3693.4]
  wire  frontend__GEN_8_4; // @[core.scala 25:25:Sodor3Stage.fir@3693.4]
  wire  frontend__GEN_11_4; // @[core.scala 25:25:Sodor3Stage.fir@3693.4]
  wire  cpath_metaReset; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath_clock; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath_io_imem_req_valid; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath_io_imem_resp_valid; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire [31:0] cpath_io_imem_resp_bits_inst; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath_io_dat_br_eq; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath_io_dat_br_lt; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath_io_dat_br_ltu; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath_io_dat_csr_eret; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath_io_ctl_exe_kill; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire [2:0] cpath_io_ctl_pc_sel; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath_io_ctl_brjmp_sel; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire [1:0] cpath_io_ctl_op1_sel; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire [1:0] cpath_io_ctl_op2_sel; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire [3:0] cpath_io_ctl_alu_fun; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire [1:0] cpath_io_ctl_wb_sel; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath_io_ctl_rf_wen; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath_io_ctl_bypassable; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire [2:0] cpath_io_ctl_csr_cmd; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath_io_ctl_dmem_fcn; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire [2:0] cpath_io_ctl_dmem_typ; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath_io_ctl_exception; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_91_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_51_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_304_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_199_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_148_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_403_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_24_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_247_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_106_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_133_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_205_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_39_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_232_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_418_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_127_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_331_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_190_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_226_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_45_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_112_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_298_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_72_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_211_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_325_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_397_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_424_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_30_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_310_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_319_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_66_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_220_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_214_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_100_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_109_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_313_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_282_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_177_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_208_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_391_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_381_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_412_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_27_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_276_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_54_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_193_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_12_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_406_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_48_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_115_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_6_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_33_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_121_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_307_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_375_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_229_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_94_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_292_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_183_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_0_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_196_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_186_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_400_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_103_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_264_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_295_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_159_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_202_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_171_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_357_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_270_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_384_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_36_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_285_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_165_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_279_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_378_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_21_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_301_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_394_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_15_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_363_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_9_3; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_258_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_97_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_345_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_339_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_18_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_147_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_330_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_86_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_273_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_351_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_231_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_189_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_153_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_288_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_366_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_252_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_180_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_71_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_174_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_168_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_372_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_3_2; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_387_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_246_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_267_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_354_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_213_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_249_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_240_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_141_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_135_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_234_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_348_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_261_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_312_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_53_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_333_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_68_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_156_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_360_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_369_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_74_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_327_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_89_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_162_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_426_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_129_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_228_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_411_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_255_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_120_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_80_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_342_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_393_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_56_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_144_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_408_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_222_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_117_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_321_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_243_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_237_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_123_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_102_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_62_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_150_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_336_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_201_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_195_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_414_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_300_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_294_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_309_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_77_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_83_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_216_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_420_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_35_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_41_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_315_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_429_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_138_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_402_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_17_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_225_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_105_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_50_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_44_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_324_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_318_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_396_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_386_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_38_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_65_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_23_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_417_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_111_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_210_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_219_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_423_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_132_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_126_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_287_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_90_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_204_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_99_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_303_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_297_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_59_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_188_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_198_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_176_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_11_3; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_380_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_93_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_161_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_192_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_207_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_405_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_260_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_26_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_114_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_269_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_182_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_399_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_368_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_390_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_32_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_281_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_275_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_291_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_47_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_5_3; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_389_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_306_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_374_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_108_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_356_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_20_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_14_2; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_29_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_82_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_170_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_185_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_278_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_143_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_96_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_263_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_164_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_158_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_362_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_377_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_257_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_284_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_179_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_383_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_242_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_8_3; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_341_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_76_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_173_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_224_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_359_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_251_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_131_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_146_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_350_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_344_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_239_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_272_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_64_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_58_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_230_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_365_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_323_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_85_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_338_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_79_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_2_3; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_245_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_70_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_152_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_167_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_422_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_371_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_266_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_125_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_212_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_254_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_155_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_149_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_227_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_113_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_140_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_326_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_425_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_404_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_353_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_248_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_107_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_311_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_73_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_67_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_347_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_206_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_410_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_419_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_233_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_305_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_128_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_332_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_88_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_52_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_46_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_134_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_221_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_407_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_382_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_28_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_40_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_55_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_329_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_194_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_392_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_236_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_101_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_61_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_34_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_116_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_122_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_320_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_215_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_335_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_293_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_428_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_49_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_137_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_200_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_209_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_95_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_413_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_314_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_308_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_16_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_395_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_385_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_104_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_302_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_317_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_203_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_172_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_197_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_370_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_416_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_22_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_271_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_119_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_379_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_187_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_401_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_43_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_296_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_286_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_364_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_1_5; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_98_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_37_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_110_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_218_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_25_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_181_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_175_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_289_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_352_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_31_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_274_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_160_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_169_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_191_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_373_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_19_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_367_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_268_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_290_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_280_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_154_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_87_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_299_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_10_4; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_398_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_4_4; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_388_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_253_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_92_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_346_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_334_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_340_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_13_3; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_256_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_328_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_81_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_355_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_7_6; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_277_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_69_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_157_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_235_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_184_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_60_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_283_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_142_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_178_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_241_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_361_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_136_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_75_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_163_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_349_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_427_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_376_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_262_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_166_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_358_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_42_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_265_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_316_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_130_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_124_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_343_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_223_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_238_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_118_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_151_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_145_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_337_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_244_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_409_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_322_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_78_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_217_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_421_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_415_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_63_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_57_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_250_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_259_1; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_139_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  cpath__GEN_84_0; // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
  wire  dpath_metaReset; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath_clock; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath_reset; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire [31:0] dpath_io_imem_req_bits_pc; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath_io_imem_resp_ready; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath_io_imem_resp_valid; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire [31:0] dpath_io_imem_resp_bits_pc; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire [31:0] dpath_io_imem_resp_bits_inst; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire [31:0] dpath_io_dmem_req_bits_addr; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire [31:0] dpath_io_dmem_req_bits_data; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath_io_dmem_req_bits_fcn; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire [2:0] dpath_io_dmem_req_bits_typ; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire [31:0] dpath_io_dmem_resp_bits_data; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath_io_ctl_exe_kill; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire [2:0] dpath_io_ctl_pc_sel; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath_io_ctl_brjmp_sel; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire [1:0] dpath_io_ctl_op1_sel; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire [1:0] dpath_io_ctl_op2_sel; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire [3:0] dpath_io_ctl_alu_fun; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire [1:0] dpath_io_ctl_wb_sel; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath_io_ctl_rf_wen; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath_io_ctl_bypassable; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire [2:0] dpath_io_ctl_csr_cmd; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath_io_ctl_dmem_fcn; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire [2:0] dpath_io_ctl_dmem_typ; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath_io_ctl_exception; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath_io_dat_br_eq; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath_io_dat_br_lt; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath_io_dat_br_ltu; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath_io_dat_csr_eret; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_338; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_224; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_218; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_21_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_323; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_302; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_6_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_239; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_317; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_385; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_197; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_12_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_296; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_9_1; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_203; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_0_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_9_2; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_212; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_320; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_200; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_388; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_191; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_181; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_190_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_15_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_289; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_299; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_311; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_206; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_367; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_175; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_305; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_274; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_373; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_376; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_382; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_370; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_349; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_262; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_355; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_277; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_194; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_184; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_293; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_157; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_3_1; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_361; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_256; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_283; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_163; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_178; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_8_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_11_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_259; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_358; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_172; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_271; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_265; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_280; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_160; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_343; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_379; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_238; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_337; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_364; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_244; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_166; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_286; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_151; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_187; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_319_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_268; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_226_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_147_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_352; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_247_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_325_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_2_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_169; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_232_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_331_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_346; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_154; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_340; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_253; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_211_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_220_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_229_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_292_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_307_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_193_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_17_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_11_2; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_313_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_328; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_2_1; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_235; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_3_3; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_23_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_250; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_208_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_214_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_241; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_5_1; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_334; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_217; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_316; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_180_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_384_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_301_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_196_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_186_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_295_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_20_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_223; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_322; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_5_2; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_279_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_310_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_285_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_202_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_378_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_351_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_387_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_189_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_14_1; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_372_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_267_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_174_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_205_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_273_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_168_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_199_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_298_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_304_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_366_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_8_2; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_360_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_288_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_375_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_255_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_261_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_270_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_150_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_333_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_177_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_381_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_1_2; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_276_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_10_1; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_354_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_348_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_249_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_369_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_183_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_282_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_162_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_156_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_165_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_7_2; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_342_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_264_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_159_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_222_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_363_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_357_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_321_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_7_3; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_330_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_243_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_237_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_315_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_336_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_258_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_171_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_303_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_146_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_13_1; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_225_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_7_4; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_231_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_240_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_339_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_153_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_252_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_297_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_324_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_219_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_1_4; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_246_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_318_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_345_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_204_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_213_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_228_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_281_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_4_2; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_0_3; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_234_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_10_3; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_312_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_192_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_306_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_207_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_16_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_22_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_300_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_327_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_182_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_291_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_290; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_4_3; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_383_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_195_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_185_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_179_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_216_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_278_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_201_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_210_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_263_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_309_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_164_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_362_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_19_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_377_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_294_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_284_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_371_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_260_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_266_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_380_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_365_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_251_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_15_2; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_359_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_152_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_188_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_173_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_287_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_386_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_245_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_272_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_344_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_198_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_167_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_254_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_3_5; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_161_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_347_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_170_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_275_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_269_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_155_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_368_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_233_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_227_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_326_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_149_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_353_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_248_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_374_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_332_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_176_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_314_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_308_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_341_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_5_5; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_18_1; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_356_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_158_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_209_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_221_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_236_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_335_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_329_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_230_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_242_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_257_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_6_5; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_350_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  wire  dpath__GEN_215_0; // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
  FrontEnd frontend ( // @[core.scala 25:25:Sodor3Stage.fir@3693.4]
    .metaReset(frontend_metaReset),
    .clock(frontend_clock),
    .reset(frontend_reset),
    .io_cpu_req_valid(frontend_io_cpu_req_valid),
    .io_cpu_req_bits_pc(frontend_io_cpu_req_bits_pc),
    .io_cpu_resp_ready(frontend_io_cpu_resp_ready),
    .io_cpu_resp_valid(frontend_io_cpu_resp_valid),
    .io_cpu_resp_bits_pc(frontend_io_cpu_resp_bits_pc),
    .io_cpu_resp_bits_inst(frontend_io_cpu_resp_bits_inst),
    .io_imem_req_bits_addr(frontend_io_imem_req_bits_addr),
    .io_imem_resp_bits_data(frontend_io_imem_resp_bits_data),
    ._GEN_1_0(frontend__GEN_1_0),
    ._GEN_10_0(frontend__GEN_10_0),
    ._GEN_13_0(frontend__GEN_13_0),
    ._GEN_7_1(frontend__GEN_7_1),
    ._GEN_9_4(frontend__GEN_9_4),
    ._GEN_12_2(frontend__GEN_12_2),
    ._GEN_6_4(frontend__GEN_6_4),
    ._GEN_14_3(frontend__GEN_14_3),
    ._GEN_5_4(frontend__GEN_5_4),
    ._GEN_8_4(frontend__GEN_8_4),
    ._GEN_11_4(frontend__GEN_11_4)
  );
  CtlPath cpath ( // @[core.scala 26:23:Sodor3Stage.fir@3696.4]
    .metaReset(cpath_metaReset),
    .clock(cpath_clock),
    .io_imem_req_valid(cpath_io_imem_req_valid),
    .io_imem_resp_valid(cpath_io_imem_resp_valid),
    .io_imem_resp_bits_inst(cpath_io_imem_resp_bits_inst),
    .io_dat_br_eq(cpath_io_dat_br_eq),
    .io_dat_br_lt(cpath_io_dat_br_lt),
    .io_dat_br_ltu(cpath_io_dat_br_ltu),
    .io_dat_csr_eret(cpath_io_dat_csr_eret),
    .io_ctl_exe_kill(cpath_io_ctl_exe_kill),
    .io_ctl_pc_sel(cpath_io_ctl_pc_sel),
    .io_ctl_brjmp_sel(cpath_io_ctl_brjmp_sel),
    .io_ctl_op1_sel(cpath_io_ctl_op1_sel),
    .io_ctl_op2_sel(cpath_io_ctl_op2_sel),
    .io_ctl_alu_fun(cpath_io_ctl_alu_fun),
    .io_ctl_wb_sel(cpath_io_ctl_wb_sel),
    .io_ctl_rf_wen(cpath_io_ctl_rf_wen),
    .io_ctl_bypassable(cpath_io_ctl_bypassable),
    .io_ctl_csr_cmd(cpath_io_ctl_csr_cmd),
    .io_ctl_dmem_fcn(cpath_io_ctl_dmem_fcn),
    .io_ctl_dmem_typ(cpath_io_ctl_dmem_typ),
    .io_ctl_exception(cpath_io_ctl_exception),
    ._GEN_91_0(cpath__GEN_91_0),
    ._GEN_51_0(cpath__GEN_51_0),
    ._GEN_304_0(cpath__GEN_304_0),
    ._GEN_199_0(cpath__GEN_199_0),
    ._GEN_148_0(cpath__GEN_148_0),
    ._GEN_403_0(cpath__GEN_403_0),
    ._GEN_24_0(cpath__GEN_24_0),
    ._GEN_247_0(cpath__GEN_247_0),
    ._GEN_106_0(cpath__GEN_106_0),
    ._GEN_133_0(cpath__GEN_133_0),
    ._GEN_205_0(cpath__GEN_205_0),
    ._GEN_39_0(cpath__GEN_39_0),
    ._GEN_232_0(cpath__GEN_232_0),
    ._GEN_418_0(cpath__GEN_418_0),
    ._GEN_127_0(cpath__GEN_127_0),
    ._GEN_331_0(cpath__GEN_331_0),
    ._GEN_190_0(cpath__GEN_190_0),
    ._GEN_226_0(cpath__GEN_226_0),
    ._GEN_45_0(cpath__GEN_45_0),
    ._GEN_112_0(cpath__GEN_112_0),
    ._GEN_298_0(cpath__GEN_298_0),
    ._GEN_72_0(cpath__GEN_72_0),
    ._GEN_211_0(cpath__GEN_211_0),
    ._GEN_325_0(cpath__GEN_325_0),
    ._GEN_397_0(cpath__GEN_397_0),
    ._GEN_424_0(cpath__GEN_424_0),
    ._GEN_30_0(cpath__GEN_30_0),
    ._GEN_310_0(cpath__GEN_310_0),
    ._GEN_319_0(cpath__GEN_319_0),
    ._GEN_66_0(cpath__GEN_66_0),
    ._GEN_220_0(cpath__GEN_220_0),
    ._GEN_214_0(cpath__GEN_214_0),
    ._GEN_100_0(cpath__GEN_100_0),
    ._GEN_109_0(cpath__GEN_109_0),
    ._GEN_313_0(cpath__GEN_313_0),
    ._GEN_282_0(cpath__GEN_282_0),
    ._GEN_177_0(cpath__GEN_177_0),
    ._GEN_208_0(cpath__GEN_208_0),
    ._GEN_391_0(cpath__GEN_391_0),
    ._GEN_381_0(cpath__GEN_381_0),
    ._GEN_412_0(cpath__GEN_412_0),
    ._GEN_27_0(cpath__GEN_27_0),
    ._GEN_276_0(cpath__GEN_276_0),
    ._GEN_54_0(cpath__GEN_54_0),
    ._GEN_193_0(cpath__GEN_193_0),
    ._GEN_12_1(cpath__GEN_12_1),
    ._GEN_406_0(cpath__GEN_406_0),
    ._GEN_48_0(cpath__GEN_48_0),
    ._GEN_115_0(cpath__GEN_115_0),
    ._GEN_6_1(cpath__GEN_6_1),
    ._GEN_33_0(cpath__GEN_33_0),
    ._GEN_121_0(cpath__GEN_121_0),
    ._GEN_307_0(cpath__GEN_307_0),
    ._GEN_375_0(cpath__GEN_375_0),
    ._GEN_229_0(cpath__GEN_229_0),
    ._GEN_94_0(cpath__GEN_94_0),
    ._GEN_292_0(cpath__GEN_292_0),
    ._GEN_183_0(cpath__GEN_183_0),
    ._GEN_0_1(cpath__GEN_0_1),
    ._GEN_196_0(cpath__GEN_196_0),
    ._GEN_186_0(cpath__GEN_186_0),
    ._GEN_400_0(cpath__GEN_400_0),
    ._GEN_103_0(cpath__GEN_103_0),
    ._GEN_264_0(cpath__GEN_264_0),
    ._GEN_295_0(cpath__GEN_295_0),
    ._GEN_159_0(cpath__GEN_159_0),
    ._GEN_202_0(cpath__GEN_202_0),
    ._GEN_171_0(cpath__GEN_171_0),
    ._GEN_357_0(cpath__GEN_357_0),
    ._GEN_270_0(cpath__GEN_270_0),
    ._GEN_384_0(cpath__GEN_384_0),
    ._GEN_36_0(cpath__GEN_36_0),
    ._GEN_285_0(cpath__GEN_285_0),
    ._GEN_165_0(cpath__GEN_165_0),
    ._GEN_279_0(cpath__GEN_279_0),
    ._GEN_378_0(cpath__GEN_378_0),
    ._GEN_21_1(cpath__GEN_21_1),
    ._GEN_301_0(cpath__GEN_301_0),
    ._GEN_394_0(cpath__GEN_394_0),
    ._GEN_15_1(cpath__GEN_15_1),
    ._GEN_363_0(cpath__GEN_363_0),
    ._GEN_9_3(cpath__GEN_9_3),
    ._GEN_258_0(cpath__GEN_258_0),
    ._GEN_97_0(cpath__GEN_97_0),
    ._GEN_345_0(cpath__GEN_345_0),
    ._GEN_339_0(cpath__GEN_339_0),
    ._GEN_18_0(cpath__GEN_18_0),
    ._GEN_147_0(cpath__GEN_147_0),
    ._GEN_330_0(cpath__GEN_330_0),
    ._GEN_86_0(cpath__GEN_86_0),
    ._GEN_273_0(cpath__GEN_273_0),
    ._GEN_351_0(cpath__GEN_351_0),
    ._GEN_231_0(cpath__GEN_231_0),
    ._GEN_189_0(cpath__GEN_189_0),
    ._GEN_153_0(cpath__GEN_153_0),
    ._GEN_288_0(cpath__GEN_288_0),
    ._GEN_366_0(cpath__GEN_366_0),
    ._GEN_252_0(cpath__GEN_252_0),
    ._GEN_180_0(cpath__GEN_180_0),
    ._GEN_71_0(cpath__GEN_71_0),
    ._GEN_174_0(cpath__GEN_174_0),
    ._GEN_168_0(cpath__GEN_168_0),
    ._GEN_372_0(cpath__GEN_372_0),
    ._GEN_3_2(cpath__GEN_3_2),
    ._GEN_387_0(cpath__GEN_387_0),
    ._GEN_246_0(cpath__GEN_246_0),
    ._GEN_267_0(cpath__GEN_267_0),
    ._GEN_354_0(cpath__GEN_354_0),
    ._GEN_213_0(cpath__GEN_213_0),
    ._GEN_249_0(cpath__GEN_249_0),
    ._GEN_240_0(cpath__GEN_240_0),
    ._GEN_141_0(cpath__GEN_141_0),
    ._GEN_135_0(cpath__GEN_135_0),
    ._GEN_234_0(cpath__GEN_234_0),
    ._GEN_348_0(cpath__GEN_348_0),
    ._GEN_261_0(cpath__GEN_261_0),
    ._GEN_312_0(cpath__GEN_312_0),
    ._GEN_53_0(cpath__GEN_53_0),
    ._GEN_333_0(cpath__GEN_333_0),
    ._GEN_68_0(cpath__GEN_68_0),
    ._GEN_156_0(cpath__GEN_156_0),
    ._GEN_360_0(cpath__GEN_360_0),
    ._GEN_369_0(cpath__GEN_369_0),
    ._GEN_74_0(cpath__GEN_74_0),
    ._GEN_327_0(cpath__GEN_327_0),
    ._GEN_89_0(cpath__GEN_89_0),
    ._GEN_162_0(cpath__GEN_162_0),
    ._GEN_426_0(cpath__GEN_426_0),
    ._GEN_129_0(cpath__GEN_129_0),
    ._GEN_228_0(cpath__GEN_228_0),
    ._GEN_411_0(cpath__GEN_411_0),
    ._GEN_255_0(cpath__GEN_255_0),
    ._GEN_120_0(cpath__GEN_120_0),
    ._GEN_80_0(cpath__GEN_80_0),
    ._GEN_342_0(cpath__GEN_342_0),
    ._GEN_393_0(cpath__GEN_393_0),
    ._GEN_56_0(cpath__GEN_56_0),
    ._GEN_144_0(cpath__GEN_144_0),
    ._GEN_408_0(cpath__GEN_408_0),
    ._GEN_222_0(cpath__GEN_222_0),
    ._GEN_117_0(cpath__GEN_117_0),
    ._GEN_321_0(cpath__GEN_321_0),
    ._GEN_243_0(cpath__GEN_243_0),
    ._GEN_237_0(cpath__GEN_237_0),
    ._GEN_123_0(cpath__GEN_123_0),
    ._GEN_102_0(cpath__GEN_102_0),
    ._GEN_62_0(cpath__GEN_62_0),
    ._GEN_150_0(cpath__GEN_150_0),
    ._GEN_336_0(cpath__GEN_336_0),
    ._GEN_201_0(cpath__GEN_201_0),
    ._GEN_195_0(cpath__GEN_195_0),
    ._GEN_414_0(cpath__GEN_414_0),
    ._GEN_300_0(cpath__GEN_300_0),
    ._GEN_294_0(cpath__GEN_294_0),
    ._GEN_309_0(cpath__GEN_309_0),
    ._GEN_77_0(cpath__GEN_77_0),
    ._GEN_83_0(cpath__GEN_83_0),
    ._GEN_216_0(cpath__GEN_216_0),
    ._GEN_420_0(cpath__GEN_420_0),
    ._GEN_35_0(cpath__GEN_35_0),
    ._GEN_41_0(cpath__GEN_41_0),
    ._GEN_315_0(cpath__GEN_315_0),
    ._GEN_429_0(cpath__GEN_429_0),
    ._GEN_138_0(cpath__GEN_138_0),
    ._GEN_402_0(cpath__GEN_402_0),
    ._GEN_17_1(cpath__GEN_17_1),
    ._GEN_225_0(cpath__GEN_225_0),
    ._GEN_105_0(cpath__GEN_105_0),
    ._GEN_50_0(cpath__GEN_50_0),
    ._GEN_44_0(cpath__GEN_44_0),
    ._GEN_324_0(cpath__GEN_324_0),
    ._GEN_318_0(cpath__GEN_318_0),
    ._GEN_396_0(cpath__GEN_396_0),
    ._GEN_386_0(cpath__GEN_386_0),
    ._GEN_38_0(cpath__GEN_38_0),
    ._GEN_65_0(cpath__GEN_65_0),
    ._GEN_23_1(cpath__GEN_23_1),
    ._GEN_417_0(cpath__GEN_417_0),
    ._GEN_111_0(cpath__GEN_111_0),
    ._GEN_210_0(cpath__GEN_210_0),
    ._GEN_219_0(cpath__GEN_219_0),
    ._GEN_423_0(cpath__GEN_423_0),
    ._GEN_132_0(cpath__GEN_132_0),
    ._GEN_126_0(cpath__GEN_126_0),
    ._GEN_287_0(cpath__GEN_287_0),
    ._GEN_90_0(cpath__GEN_90_0),
    ._GEN_204_0(cpath__GEN_204_0),
    ._GEN_99_0(cpath__GEN_99_0),
    ._GEN_303_0(cpath__GEN_303_0),
    ._GEN_297_0(cpath__GEN_297_0),
    ._GEN_59_0(cpath__GEN_59_0),
    ._GEN_188_0(cpath__GEN_188_0),
    ._GEN_198_0(cpath__GEN_198_0),
    ._GEN_176_0(cpath__GEN_176_0),
    ._GEN_11_3(cpath__GEN_11_3),
    ._GEN_380_0(cpath__GEN_380_0),
    ._GEN_93_0(cpath__GEN_93_0),
    ._GEN_161_0(cpath__GEN_161_0),
    ._GEN_192_0(cpath__GEN_192_0),
    ._GEN_207_0(cpath__GEN_207_0),
    ._GEN_405_0(cpath__GEN_405_0),
    ._GEN_260_0(cpath__GEN_260_0),
    ._GEN_26_0(cpath__GEN_26_0),
    ._GEN_114_0(cpath__GEN_114_0),
    ._GEN_269_0(cpath__GEN_269_0),
    ._GEN_182_0(cpath__GEN_182_0),
    ._GEN_399_0(cpath__GEN_399_0),
    ._GEN_368_0(cpath__GEN_368_0),
    ._GEN_390_0(cpath__GEN_390_0),
    ._GEN_32_0(cpath__GEN_32_0),
    ._GEN_281_0(cpath__GEN_281_0),
    ._GEN_275_0(cpath__GEN_275_0),
    ._GEN_291_0(cpath__GEN_291_0),
    ._GEN_47_0(cpath__GEN_47_0),
    ._GEN_5_3(cpath__GEN_5_3),
    ._GEN_389_0(cpath__GEN_389_0),
    ._GEN_306_0(cpath__GEN_306_0),
    ._GEN_374_0(cpath__GEN_374_0),
    ._GEN_108_0(cpath__GEN_108_0),
    ._GEN_356_0(cpath__GEN_356_0),
    ._GEN_20_1(cpath__GEN_20_1),
    ._GEN_14_2(cpath__GEN_14_2),
    ._GEN_29_0(cpath__GEN_29_0),
    ._GEN_82_0(cpath__GEN_82_0),
    ._GEN_170_0(cpath__GEN_170_0),
    ._GEN_185_0(cpath__GEN_185_0),
    ._GEN_278_0(cpath__GEN_278_0),
    ._GEN_143_0(cpath__GEN_143_0),
    ._GEN_96_0(cpath__GEN_96_0),
    ._GEN_263_0(cpath__GEN_263_0),
    ._GEN_164_0(cpath__GEN_164_0),
    ._GEN_158_0(cpath__GEN_158_0),
    ._GEN_362_0(cpath__GEN_362_0),
    ._GEN_377_0(cpath__GEN_377_0),
    ._GEN_257_0(cpath__GEN_257_0),
    ._GEN_284_0(cpath__GEN_284_0),
    ._GEN_179_0(cpath__GEN_179_0),
    ._GEN_383_0(cpath__GEN_383_0),
    ._GEN_242_0(cpath__GEN_242_0),
    ._GEN_8_3(cpath__GEN_8_3),
    ._GEN_341_0(cpath__GEN_341_0),
    ._GEN_76_0(cpath__GEN_76_0),
    ._GEN_173_0(cpath__GEN_173_0),
    ._GEN_224_1(cpath__GEN_224_1),
    ._GEN_359_0(cpath__GEN_359_0),
    ._GEN_251_0(cpath__GEN_251_0),
    ._GEN_131_0(cpath__GEN_131_0),
    ._GEN_146_0(cpath__GEN_146_0),
    ._GEN_350_0(cpath__GEN_350_0),
    ._GEN_344_0(cpath__GEN_344_0),
    ._GEN_239_1(cpath__GEN_239_1),
    ._GEN_272_0(cpath__GEN_272_0),
    ._GEN_64_0(cpath__GEN_64_0),
    ._GEN_58_0(cpath__GEN_58_0),
    ._GEN_230_0(cpath__GEN_230_0),
    ._GEN_365_0(cpath__GEN_365_0),
    ._GEN_323_1(cpath__GEN_323_1),
    ._GEN_85_0(cpath__GEN_85_0),
    ._GEN_338_1(cpath__GEN_338_1),
    ._GEN_79_0(cpath__GEN_79_0),
    ._GEN_2_3(cpath__GEN_2_3),
    ._GEN_245_0(cpath__GEN_245_0),
    ._GEN_70_0(cpath__GEN_70_0),
    ._GEN_152_0(cpath__GEN_152_0),
    ._GEN_167_0(cpath__GEN_167_0),
    ._GEN_422_0(cpath__GEN_422_0),
    ._GEN_371_0(cpath__GEN_371_0),
    ._GEN_266_0(cpath__GEN_266_0),
    ._GEN_125_0(cpath__GEN_125_0),
    ._GEN_212_1(cpath__GEN_212_1),
    ._GEN_254_0(cpath__GEN_254_0),
    ._GEN_155_0(cpath__GEN_155_0),
    ._GEN_149_0(cpath__GEN_149_0),
    ._GEN_227_0(cpath__GEN_227_0),
    ._GEN_113_0(cpath__GEN_113_0),
    ._GEN_140_0(cpath__GEN_140_0),
    ._GEN_326_0(cpath__GEN_326_0),
    ._GEN_425_0(cpath__GEN_425_0),
    ._GEN_404_0(cpath__GEN_404_0),
    ._GEN_353_0(cpath__GEN_353_0),
    ._GEN_248_0(cpath__GEN_248_0),
    ._GEN_107_0(cpath__GEN_107_0),
    ._GEN_311_1(cpath__GEN_311_1),
    ._GEN_73_0(cpath__GEN_73_0),
    ._GEN_67_0(cpath__GEN_67_0),
    ._GEN_347_0(cpath__GEN_347_0),
    ._GEN_206_1(cpath__GEN_206_1),
    ._GEN_410_0(cpath__GEN_410_0),
    ._GEN_419_0(cpath__GEN_419_0),
    ._GEN_233_0(cpath__GEN_233_0),
    ._GEN_305_1(cpath__GEN_305_1),
    ._GEN_128_0(cpath__GEN_128_0),
    ._GEN_332_0(cpath__GEN_332_0),
    ._GEN_88_0(cpath__GEN_88_0),
    ._GEN_52_0(cpath__GEN_52_0),
    ._GEN_46_0(cpath__GEN_46_0),
    ._GEN_134_0(cpath__GEN_134_0),
    ._GEN_221_0(cpath__GEN_221_0),
    ._GEN_407_0(cpath__GEN_407_0),
    ._GEN_382_1(cpath__GEN_382_1),
    ._GEN_28_0(cpath__GEN_28_0),
    ._GEN_40_0(cpath__GEN_40_0),
    ._GEN_55_0(cpath__GEN_55_0),
    ._GEN_329_0(cpath__GEN_329_0),
    ._GEN_194_1(cpath__GEN_194_1),
    ._GEN_392_0(cpath__GEN_392_0),
    ._GEN_236_0(cpath__GEN_236_0),
    ._GEN_101_0(cpath__GEN_101_0),
    ._GEN_61_0(cpath__GEN_61_0),
    ._GEN_34_0(cpath__GEN_34_0),
    ._GEN_116_0(cpath__GEN_116_0),
    ._GEN_122_0(cpath__GEN_122_0),
    ._GEN_320_1(cpath__GEN_320_1),
    ._GEN_215_0(cpath__GEN_215_0),
    ._GEN_335_0(cpath__GEN_335_0),
    ._GEN_293_1(cpath__GEN_293_1),
    ._GEN_428_0(cpath__GEN_428_0),
    ._GEN_49_0(cpath__GEN_49_0),
    ._GEN_137_0(cpath__GEN_137_0),
    ._GEN_200_1(cpath__GEN_200_1),
    ._GEN_209_0(cpath__GEN_209_0),
    ._GEN_95_0(cpath__GEN_95_0),
    ._GEN_413_0(cpath__GEN_413_0),
    ._GEN_314_0(cpath__GEN_314_0),
    ._GEN_308_0(cpath__GEN_308_0),
    ._GEN_16_1(cpath__GEN_16_1),
    ._GEN_395_0(cpath__GEN_395_0),
    ._GEN_385_1(cpath__GEN_385_1),
    ._GEN_104_0(cpath__GEN_104_0),
    ._GEN_302_1(cpath__GEN_302_1),
    ._GEN_317_1(cpath__GEN_317_1),
    ._GEN_203_1(cpath__GEN_203_1),
    ._GEN_172_1(cpath__GEN_172_1),
    ._GEN_197_1(cpath__GEN_197_1),
    ._GEN_370_1(cpath__GEN_370_1),
    ._GEN_416_0(cpath__GEN_416_0),
    ._GEN_22_1(cpath__GEN_22_1),
    ._GEN_271_1(cpath__GEN_271_1),
    ._GEN_119_0(cpath__GEN_119_0),
    ._GEN_379_1(cpath__GEN_379_1),
    ._GEN_187_1(cpath__GEN_187_1),
    ._GEN_401_0(cpath__GEN_401_0),
    ._GEN_43_0(cpath__GEN_43_0),
    ._GEN_296_1(cpath__GEN_296_1),
    ._GEN_286_1(cpath__GEN_286_1),
    ._GEN_364_1(cpath__GEN_364_1),
    ._GEN_1_5(cpath__GEN_1_5),
    ._GEN_98_0(cpath__GEN_98_0),
    ._GEN_37_0(cpath__GEN_37_0),
    ._GEN_110_0(cpath__GEN_110_0),
    ._GEN_218_1(cpath__GEN_218_1),
    ._GEN_25_0(cpath__GEN_25_0),
    ._GEN_181_1(cpath__GEN_181_1),
    ._GEN_175_1(cpath__GEN_175_1),
    ._GEN_289_1(cpath__GEN_289_1),
    ._GEN_352_1(cpath__GEN_352_1),
    ._GEN_31_0(cpath__GEN_31_0),
    ._GEN_274_1(cpath__GEN_274_1),
    ._GEN_160_1(cpath__GEN_160_1),
    ._GEN_169_1(cpath__GEN_169_1),
    ._GEN_191_1(cpath__GEN_191_1),
    ._GEN_373_1(cpath__GEN_373_1),
    ._GEN_19_1(cpath__GEN_19_1),
    ._GEN_367_1(cpath__GEN_367_1),
    ._GEN_268_1(cpath__GEN_268_1),
    ._GEN_290_1(cpath__GEN_290_1),
    ._GEN_280_1(cpath__GEN_280_1),
    ._GEN_154_1(cpath__GEN_154_1),
    ._GEN_87_0(cpath__GEN_87_0),
    ._GEN_299_1(cpath__GEN_299_1),
    ._GEN_10_4(cpath__GEN_10_4),
    ._GEN_398_0(cpath__GEN_398_0),
    ._GEN_4_4(cpath__GEN_4_4),
    ._GEN_388_1(cpath__GEN_388_1),
    ._GEN_253_1(cpath__GEN_253_1),
    ._GEN_92_0(cpath__GEN_92_0),
    ._GEN_346_1(cpath__GEN_346_1),
    ._GEN_334_1(cpath__GEN_334_1),
    ._GEN_340_1(cpath__GEN_340_1),
    ._GEN_13_3(cpath__GEN_13_3),
    ._GEN_256_1(cpath__GEN_256_1),
    ._GEN_328_1(cpath__GEN_328_1),
    ._GEN_81_0(cpath__GEN_81_0),
    ._GEN_355_1(cpath__GEN_355_1),
    ._GEN_7_6(cpath__GEN_7_6),
    ._GEN_277_1(cpath__GEN_277_1),
    ._GEN_69_0(cpath__GEN_69_0),
    ._GEN_157_1(cpath__GEN_157_1),
    ._GEN_235_1(cpath__GEN_235_1),
    ._GEN_184_1(cpath__GEN_184_1),
    ._GEN_60_0(cpath__GEN_60_0),
    ._GEN_283_1(cpath__GEN_283_1),
    ._GEN_142_0(cpath__GEN_142_0),
    ._GEN_178_1(cpath__GEN_178_1),
    ._GEN_241_1(cpath__GEN_241_1),
    ._GEN_361_1(cpath__GEN_361_1),
    ._GEN_136_0(cpath__GEN_136_0),
    ._GEN_75_0(cpath__GEN_75_0),
    ._GEN_163_1(cpath__GEN_163_1),
    ._GEN_349_1(cpath__GEN_349_1),
    ._GEN_427_0(cpath__GEN_427_0),
    ._GEN_376_1(cpath__GEN_376_1),
    ._GEN_262_1(cpath__GEN_262_1),
    ._GEN_166_1(cpath__GEN_166_1),
    ._GEN_358_1(cpath__GEN_358_1),
    ._GEN_42_0(cpath__GEN_42_0),
    ._GEN_265_1(cpath__GEN_265_1),
    ._GEN_316_1(cpath__GEN_316_1),
    ._GEN_130_0(cpath__GEN_130_0),
    ._GEN_124_0(cpath__GEN_124_0),
    ._GEN_343_1(cpath__GEN_343_1),
    ._GEN_223_1(cpath__GEN_223_1),
    ._GEN_238_1(cpath__GEN_238_1),
    ._GEN_118_0(cpath__GEN_118_0),
    ._GEN_151_1(cpath__GEN_151_1),
    ._GEN_145_0(cpath__GEN_145_0),
    ._GEN_337_1(cpath__GEN_337_1),
    ._GEN_244_1(cpath__GEN_244_1),
    ._GEN_409_0(cpath__GEN_409_0),
    ._GEN_322_1(cpath__GEN_322_1),
    ._GEN_78_0(cpath__GEN_78_0),
    ._GEN_217_1(cpath__GEN_217_1),
    ._GEN_421_0(cpath__GEN_421_0),
    ._GEN_415_0(cpath__GEN_415_0),
    ._GEN_63_0(cpath__GEN_63_0),
    ._GEN_57_0(cpath__GEN_57_0),
    ._GEN_250_1(cpath__GEN_250_1),
    ._GEN_259_1(cpath__GEN_259_1),
    ._GEN_139_0(cpath__GEN_139_0),
    ._GEN_84_0(cpath__GEN_84_0)
  );
  DatPath dpath ( // @[core.scala 27:23:Sodor3Stage.fir@3699.4]
    .metaReset(dpath_metaReset),
    .clock(dpath_clock),
    .reset(dpath_reset),
    .io_imem_req_bits_pc(dpath_io_imem_req_bits_pc),
    .io_imem_resp_ready(dpath_io_imem_resp_ready),
    .io_imem_resp_valid(dpath_io_imem_resp_valid),
    .io_imem_resp_bits_pc(dpath_io_imem_resp_bits_pc),
    .io_imem_resp_bits_inst(dpath_io_imem_resp_bits_inst),
    .io_dmem_req_bits_addr(dpath_io_dmem_req_bits_addr),
    .io_dmem_req_bits_data(dpath_io_dmem_req_bits_data),
    .io_dmem_req_bits_fcn(dpath_io_dmem_req_bits_fcn),
    .io_dmem_req_bits_typ(dpath_io_dmem_req_bits_typ),
    .io_dmem_resp_bits_data(dpath_io_dmem_resp_bits_data),
    .io_ctl_exe_kill(dpath_io_ctl_exe_kill),
    .io_ctl_pc_sel(dpath_io_ctl_pc_sel),
    .io_ctl_brjmp_sel(dpath_io_ctl_brjmp_sel),
    .io_ctl_op1_sel(dpath_io_ctl_op1_sel),
    .io_ctl_op2_sel(dpath_io_ctl_op2_sel),
    .io_ctl_alu_fun(dpath_io_ctl_alu_fun),
    .io_ctl_wb_sel(dpath_io_ctl_wb_sel),
    .io_ctl_rf_wen(dpath_io_ctl_rf_wen),
    .io_ctl_bypassable(dpath_io_ctl_bypassable),
    .io_ctl_csr_cmd(dpath_io_ctl_csr_cmd),
    .io_ctl_dmem_fcn(dpath_io_ctl_dmem_fcn),
    .io_ctl_dmem_typ(dpath_io_ctl_dmem_typ),
    .io_ctl_exception(dpath_io_ctl_exception),
    .io_dat_br_eq(dpath_io_dat_br_eq),
    .io_dat_br_lt(dpath_io_dat_br_lt),
    .io_dat_br_ltu(dpath_io_dat_br_ltu),
    .io_dat_csr_eret(dpath_io_dat_csr_eret),
    ._GEN_338(dpath__GEN_338),
    ._GEN_224(dpath__GEN_224),
    ._GEN_218(dpath__GEN_218),
    ._GEN_21_0(dpath__GEN_21_0),
    ._GEN_323(dpath__GEN_323),
    ._GEN_302(dpath__GEN_302),
    ._GEN_6_0(dpath__GEN_6_0),
    ._GEN_239(dpath__GEN_239),
    ._GEN_317(dpath__GEN_317),
    ._GEN_385(dpath__GEN_385),
    ._GEN_197(dpath__GEN_197),
    ._GEN_12_0(dpath__GEN_12_0),
    ._GEN_296(dpath__GEN_296),
    ._GEN_9_1(dpath__GEN_9_1),
    ._GEN_203(dpath__GEN_203),
    ._GEN_0_0(dpath__GEN_0_0),
    ._GEN_9_2(dpath__GEN_9_2),
    ._GEN_212(dpath__GEN_212),
    ._GEN_320(dpath__GEN_320),
    ._GEN_200(dpath__GEN_200),
    ._GEN_388(dpath__GEN_388),
    ._GEN_191(dpath__GEN_191),
    ._GEN_181(dpath__GEN_181),
    ._GEN_190_0(dpath__GEN_190_0),
    ._GEN_15_0(dpath__GEN_15_0),
    ._GEN_289(dpath__GEN_289),
    ._GEN_299(dpath__GEN_299),
    ._GEN_311(dpath__GEN_311),
    ._GEN_206(dpath__GEN_206),
    ._GEN_367(dpath__GEN_367),
    ._GEN_175(dpath__GEN_175),
    ._GEN_305(dpath__GEN_305),
    ._GEN_274(dpath__GEN_274),
    ._GEN_373(dpath__GEN_373),
    ._GEN_376(dpath__GEN_376),
    ._GEN_382(dpath__GEN_382),
    ._GEN_370(dpath__GEN_370),
    ._GEN_349(dpath__GEN_349),
    ._GEN_262(dpath__GEN_262),
    ._GEN_355(dpath__GEN_355),
    ._GEN_277(dpath__GEN_277),
    ._GEN_194(dpath__GEN_194),
    ._GEN_184(dpath__GEN_184),
    ._GEN_293(dpath__GEN_293),
    ._GEN_157(dpath__GEN_157),
    ._GEN_3_1(dpath__GEN_3_1),
    ._GEN_361(dpath__GEN_361),
    ._GEN_256(dpath__GEN_256),
    ._GEN_283(dpath__GEN_283),
    ._GEN_163(dpath__GEN_163),
    ._GEN_178(dpath__GEN_178),
    ._GEN_8_0(dpath__GEN_8_0),
    ._GEN_11_0(dpath__GEN_11_0),
    ._GEN_259(dpath__GEN_259),
    ._GEN_358(dpath__GEN_358),
    ._GEN_172(dpath__GEN_172),
    ._GEN_271(dpath__GEN_271),
    ._GEN_265(dpath__GEN_265),
    ._GEN_280(dpath__GEN_280),
    ._GEN_160(dpath__GEN_160),
    ._GEN_343(dpath__GEN_343),
    ._GEN_379(dpath__GEN_379),
    ._GEN_238(dpath__GEN_238),
    ._GEN_337(dpath__GEN_337),
    ._GEN_364(dpath__GEN_364),
    ._GEN_244(dpath__GEN_244),
    ._GEN_166(dpath__GEN_166),
    ._GEN_286(dpath__GEN_286),
    ._GEN_151(dpath__GEN_151),
    ._GEN_187(dpath__GEN_187),
    ._GEN_319_0(dpath__GEN_319_0),
    ._GEN_268(dpath__GEN_268),
    ._GEN_226_0(dpath__GEN_226_0),
    ._GEN_147_0(dpath__GEN_147_0),
    ._GEN_352(dpath__GEN_352),
    ._GEN_247_0(dpath__GEN_247_0),
    ._GEN_325_0(dpath__GEN_325_0),
    ._GEN_2_0(dpath__GEN_2_0),
    ._GEN_169(dpath__GEN_169),
    ._GEN_232_0(dpath__GEN_232_0),
    ._GEN_331_0(dpath__GEN_331_0),
    ._GEN_346(dpath__GEN_346),
    ._GEN_154(dpath__GEN_154),
    ._GEN_340(dpath__GEN_340),
    ._GEN_253(dpath__GEN_253),
    ._GEN_211_0(dpath__GEN_211_0),
    ._GEN_220_0(dpath__GEN_220_0),
    ._GEN_229_0(dpath__GEN_229_0),
    ._GEN_292_0(dpath__GEN_292_0),
    ._GEN_307_0(dpath__GEN_307_0),
    ._GEN_193_0(dpath__GEN_193_0),
    ._GEN_17_0(dpath__GEN_17_0),
    ._GEN_11_2(dpath__GEN_11_2),
    ._GEN_313_0(dpath__GEN_313_0),
    ._GEN_328(dpath__GEN_328),
    ._GEN_2_1(dpath__GEN_2_1),
    ._GEN_235(dpath__GEN_235),
    ._GEN_3_3(dpath__GEN_3_3),
    ._GEN_23_0(dpath__GEN_23_0),
    ._GEN_250(dpath__GEN_250),
    ._GEN_208_0(dpath__GEN_208_0),
    ._GEN_214_0(dpath__GEN_214_0),
    ._GEN_241(dpath__GEN_241),
    ._GEN_5_1(dpath__GEN_5_1),
    ._GEN_334(dpath__GEN_334),
    ._GEN_217(dpath__GEN_217),
    ._GEN_316(dpath__GEN_316),
    ._GEN_180_0(dpath__GEN_180_0),
    ._GEN_384_0(dpath__GEN_384_0),
    ._GEN_301_0(dpath__GEN_301_0),
    ._GEN_196_0(dpath__GEN_196_0),
    ._GEN_186_0(dpath__GEN_186_0),
    ._GEN_295_0(dpath__GEN_295_0),
    ._GEN_20_0(dpath__GEN_20_0),
    ._GEN_223(dpath__GEN_223),
    ._GEN_322(dpath__GEN_322),
    ._GEN_5_2(dpath__GEN_5_2),
    ._GEN_279_0(dpath__GEN_279_0),
    ._GEN_310_0(dpath__GEN_310_0),
    ._GEN_285_0(dpath__GEN_285_0),
    ._GEN_202_0(dpath__GEN_202_0),
    ._GEN_378_0(dpath__GEN_378_0),
    ._GEN_351_0(dpath__GEN_351_0),
    ._GEN_387_0(dpath__GEN_387_0),
    ._GEN_189_0(dpath__GEN_189_0),
    ._GEN_14_1(dpath__GEN_14_1),
    ._GEN_372_0(dpath__GEN_372_0),
    ._GEN_267_0(dpath__GEN_267_0),
    ._GEN_174_0(dpath__GEN_174_0),
    ._GEN_205_0(dpath__GEN_205_0),
    ._GEN_273_0(dpath__GEN_273_0),
    ._GEN_168_0(dpath__GEN_168_0),
    ._GEN_199_0(dpath__GEN_199_0),
    ._GEN_298_0(dpath__GEN_298_0),
    ._GEN_304_0(dpath__GEN_304_0),
    ._GEN_366_0(dpath__GEN_366_0),
    ._GEN_8_2(dpath__GEN_8_2),
    ._GEN_360_0(dpath__GEN_360_0),
    ._GEN_288_0(dpath__GEN_288_0),
    ._GEN_375_0(dpath__GEN_375_0),
    ._GEN_255_0(dpath__GEN_255_0),
    ._GEN_261_0(dpath__GEN_261_0),
    ._GEN_270_0(dpath__GEN_270_0),
    ._GEN_150_0(dpath__GEN_150_0),
    ._GEN_333_0(dpath__GEN_333_0),
    ._GEN_177_0(dpath__GEN_177_0),
    ._GEN_381_0(dpath__GEN_381_0),
    ._GEN_1_2(dpath__GEN_1_2),
    ._GEN_276_0(dpath__GEN_276_0),
    ._GEN_10_1(dpath__GEN_10_1),
    ._GEN_354_0(dpath__GEN_354_0),
    ._GEN_348_0(dpath__GEN_348_0),
    ._GEN_249_0(dpath__GEN_249_0),
    ._GEN_369_0(dpath__GEN_369_0),
    ._GEN_183_0(dpath__GEN_183_0),
    ._GEN_282_0(dpath__GEN_282_0),
    ._GEN_162_0(dpath__GEN_162_0),
    ._GEN_156_0(dpath__GEN_156_0),
    ._GEN_165_0(dpath__GEN_165_0),
    ._GEN_7_2(dpath__GEN_7_2),
    ._GEN_342_0(dpath__GEN_342_0),
    ._GEN_264_0(dpath__GEN_264_0),
    ._GEN_159_0(dpath__GEN_159_0),
    ._GEN_222_0(dpath__GEN_222_0),
    ._GEN_363_0(dpath__GEN_363_0),
    ._GEN_357_0(dpath__GEN_357_0),
    ._GEN_321_0(dpath__GEN_321_0),
    ._GEN_7_3(dpath__GEN_7_3),
    ._GEN_330_0(dpath__GEN_330_0),
    ._GEN_243_0(dpath__GEN_243_0),
    ._GEN_237_0(dpath__GEN_237_0),
    ._GEN_315_0(dpath__GEN_315_0),
    ._GEN_336_0(dpath__GEN_336_0),
    ._GEN_258_0(dpath__GEN_258_0),
    ._GEN_171_0(dpath__GEN_171_0),
    ._GEN_303_0(dpath__GEN_303_0),
    ._GEN_146_0(dpath__GEN_146_0),
    ._GEN_13_1(dpath__GEN_13_1),
    ._GEN_225_0(dpath__GEN_225_0),
    ._GEN_7_4(dpath__GEN_7_4),
    ._GEN_231_0(dpath__GEN_231_0),
    ._GEN_240_0(dpath__GEN_240_0),
    ._GEN_339_0(dpath__GEN_339_0),
    ._GEN_153_0(dpath__GEN_153_0),
    ._GEN_252_0(dpath__GEN_252_0),
    ._GEN_297_0(dpath__GEN_297_0),
    ._GEN_324_0(dpath__GEN_324_0),
    ._GEN_219_0(dpath__GEN_219_0),
    ._GEN_1_4(dpath__GEN_1_4),
    ._GEN_246_0(dpath__GEN_246_0),
    ._GEN_318_0(dpath__GEN_318_0),
    ._GEN_345_0(dpath__GEN_345_0),
    ._GEN_204_0(dpath__GEN_204_0),
    ._GEN_213_0(dpath__GEN_213_0),
    ._GEN_228_0(dpath__GEN_228_0),
    ._GEN_281_0(dpath__GEN_281_0),
    ._GEN_4_2(dpath__GEN_4_2),
    ._GEN_0_3(dpath__GEN_0_3),
    ._GEN_234_0(dpath__GEN_234_0),
    ._GEN_10_3(dpath__GEN_10_3),
    ._GEN_312_0(dpath__GEN_312_0),
    ._GEN_192_0(dpath__GEN_192_0),
    ._GEN_306_0(dpath__GEN_306_0),
    ._GEN_207_0(dpath__GEN_207_0),
    ._GEN_16_0(dpath__GEN_16_0),
    ._GEN_22_0(dpath__GEN_22_0),
    ._GEN_300_0(dpath__GEN_300_0),
    ._GEN_327_0(dpath__GEN_327_0),
    ._GEN_182_0(dpath__GEN_182_0),
    ._GEN_291_0(dpath__GEN_291_0),
    ._GEN_290(dpath__GEN_290),
    ._GEN_4_3(dpath__GEN_4_3),
    ._GEN_383_0(dpath__GEN_383_0),
    ._GEN_195_0(dpath__GEN_195_0),
    ._GEN_185_0(dpath__GEN_185_0),
    ._GEN_179_0(dpath__GEN_179_0),
    ._GEN_216_0(dpath__GEN_216_0),
    ._GEN_278_0(dpath__GEN_278_0),
    ._GEN_201_0(dpath__GEN_201_0),
    ._GEN_210_0(dpath__GEN_210_0),
    ._GEN_263_0(dpath__GEN_263_0),
    ._GEN_309_0(dpath__GEN_309_0),
    ._GEN_164_0(dpath__GEN_164_0),
    ._GEN_362_0(dpath__GEN_362_0),
    ._GEN_19_0(dpath__GEN_19_0),
    ._GEN_377_0(dpath__GEN_377_0),
    ._GEN_294_0(dpath__GEN_294_0),
    ._GEN_284_0(dpath__GEN_284_0),
    ._GEN_371_0(dpath__GEN_371_0),
    ._GEN_260_0(dpath__GEN_260_0),
    ._GEN_266_0(dpath__GEN_266_0),
    ._GEN_380_0(dpath__GEN_380_0),
    ._GEN_365_0(dpath__GEN_365_0),
    ._GEN_251_0(dpath__GEN_251_0),
    ._GEN_15_2(dpath__GEN_15_2),
    ._GEN_359_0(dpath__GEN_359_0),
    ._GEN_152_0(dpath__GEN_152_0),
    ._GEN_188_0(dpath__GEN_188_0),
    ._GEN_173_0(dpath__GEN_173_0),
    ._GEN_287_0(dpath__GEN_287_0),
    ._GEN_386_0(dpath__GEN_386_0),
    ._GEN_245_0(dpath__GEN_245_0),
    ._GEN_272_0(dpath__GEN_272_0),
    ._GEN_344_0(dpath__GEN_344_0),
    ._GEN_198_0(dpath__GEN_198_0),
    ._GEN_167_0(dpath__GEN_167_0),
    ._GEN_254_0(dpath__GEN_254_0),
    ._GEN_3_5(dpath__GEN_3_5),
    ._GEN_161_0(dpath__GEN_161_0),
    ._GEN_347_0(dpath__GEN_347_0),
    ._GEN_170_0(dpath__GEN_170_0),
    ._GEN_275_0(dpath__GEN_275_0),
    ._GEN_269_0(dpath__GEN_269_0),
    ._GEN_155_0(dpath__GEN_155_0),
    ._GEN_368_0(dpath__GEN_368_0),
    ._GEN_233_0(dpath__GEN_233_0),
    ._GEN_227_0(dpath__GEN_227_0),
    ._GEN_326_0(dpath__GEN_326_0),
    ._GEN_149_0(dpath__GEN_149_0),
    ._GEN_353_0(dpath__GEN_353_0),
    ._GEN_248_0(dpath__GEN_248_0),
    ._GEN_374_0(dpath__GEN_374_0),
    ._GEN_332_0(dpath__GEN_332_0),
    ._GEN_176_0(dpath__GEN_176_0),
    ._GEN_314_0(dpath__GEN_314_0),
    ._GEN_308_0(dpath__GEN_308_0),
    ._GEN_341_0(dpath__GEN_341_0),
    ._GEN_5_5(dpath__GEN_5_5),
    ._GEN_18_1(dpath__GEN_18_1),
    ._GEN_356_0(dpath__GEN_356_0),
    ._GEN_158_0(dpath__GEN_158_0),
    ._GEN_209_0(dpath__GEN_209_0),
    ._GEN_221_0(dpath__GEN_221_0),
    ._GEN_236_0(dpath__GEN_236_0),
    ._GEN_335_0(dpath__GEN_335_0),
    ._GEN_329_0(dpath__GEN_329_0),
    ._GEN_230_0(dpath__GEN_230_0),
    ._GEN_242_0(dpath__GEN_242_0),
    ._GEN_257_0(dpath__GEN_257_0),
    ._GEN_6_5(dpath__GEN_6_5),
    ._GEN_350_0(dpath__GEN_350_0),
    ._GEN_215_0(dpath__GEN_215_0)
  );
  assign frontend_metaReset = metaReset;
  assign cpath_metaReset = metaReset;
  assign dpath_metaReset = metaReset;
  assign io_imem_req_bits_addr = frontend_io_imem_req_bits_addr;
  assign io_dmem_req_bits_addr = dpath_io_dmem_req_bits_addr;
  assign io_dmem_req_bits_data = dpath_io_dmem_req_bits_data;
  assign io_dmem_req_bits_fcn = dpath_io_dmem_req_bits_fcn;
  assign io_dmem_req_bits_typ = dpath_io_dmem_req_bits_typ;
  assign _GEN_338 = dpath__GEN_338;
  assign _GEN_224 = dpath__GEN_224;
  assign _GEN_218 = dpath__GEN_218;
  assign _GEN_21 = dpath__GEN_21_0;
  assign _GEN_91 = cpath__GEN_91_0;
  assign _GEN_323 = dpath__GEN_323;
  assign _GEN_302 = dpath__GEN_302;
  assign _GEN_51 = cpath__GEN_51_0;
  assign _GEN_304 = cpath__GEN_304_0;
  assign _GEN_199 = cpath__GEN_199_0;
  assign _GEN_6 = dpath__GEN_6_0;
  assign _GEN_148 = cpath__GEN_148_0;
  assign _GEN_239 = dpath__GEN_239;
  assign _GEN_403 = cpath__GEN_403_0;
  assign _GEN_1 = frontend__GEN_1_0;
  assign _GEN_24 = cpath__GEN_24_0;
  assign _GEN_247 = cpath__GEN_247_0;
  assign _GEN_106 = cpath__GEN_106_0;
  assign _GEN_317 = dpath__GEN_317;
  assign _GEN_133 = cpath__GEN_133_0;
  assign _GEN_205 = cpath__GEN_205_0;
  assign _GEN_385 = dpath__GEN_385;
  assign _GEN_39 = cpath__GEN_39_0;
  assign _GEN_232 = cpath__GEN_232_0;
  assign _GEN_418 = cpath__GEN_418_0;
  assign _GEN_127 = cpath__GEN_127_0;
  assign _GEN_197 = dpath__GEN_197;
  assign _GEN_331 = cpath__GEN_331_0;
  assign _GEN_190 = cpath__GEN_190_0;
  assign _GEN_12 = dpath__GEN_12_0;
  assign _GEN_226 = cpath__GEN_226_0;
  assign _GEN_296 = dpath__GEN_296;
  assign _GEN_9_0 = dpath__GEN_9_1;
  assign _GEN_45 = cpath__GEN_45_0;
  assign _GEN_112 = cpath__GEN_112_0;
  assign _GEN_298 = cpath__GEN_298_0;
  assign _GEN_203 = dpath__GEN_203;
  assign _GEN_72 = cpath__GEN_72_0;
  assign _GEN_211 = cpath__GEN_211_0;
  assign _GEN_325 = cpath__GEN_325_0;
  assign _GEN_397 = cpath__GEN_397_0;
  assign _GEN_0 = dpath__GEN_0_0;
  assign _GEN_424 = cpath__GEN_424_0;
  assign _GEN_30 = cpath__GEN_30_0;
  assign _GEN_310 = cpath__GEN_310_0;
  assign _GEN_319 = cpath__GEN_319_0;
  assign _GEN_66 = cpath__GEN_66_0;
  assign _GEN_9_1 = dpath__GEN_9_2;
  assign _GEN_212 = dpath__GEN_212;
  assign _GEN_220 = cpath__GEN_220_0;
  assign _GEN_214 = cpath__GEN_214_0;
  assign _GEN_100 = cpath__GEN_100_0;
  assign _GEN_109 = cpath__GEN_109_0;
  assign _GEN_320 = dpath__GEN_320;
  assign _GEN_313 = cpath__GEN_313_0;
  assign _GEN_282 = cpath__GEN_282_0;
  assign _GEN_200 = dpath__GEN_200;
  assign _GEN_177 = cpath__GEN_177_0;
  assign _GEN_208 = cpath__GEN_208_0;
  assign _GEN_388 = dpath__GEN_388;
  assign _GEN_391 = cpath__GEN_391_0;
  assign _GEN_381 = cpath__GEN_381_0;
  assign _GEN_412 = cpath__GEN_412_0;
  assign _GEN_27 = cpath__GEN_27_0;
  assign _GEN_276 = cpath__GEN_276_0;
  assign _GEN_191 = dpath__GEN_191;
  assign _GEN_181 = dpath__GEN_181;
  assign _GEN_54 = cpath__GEN_54_0;
  assign _GEN_193 = cpath__GEN_193_0;
  assign _GEN_190_0 = dpath__GEN_190_0;
  assign _GEN_15 = dpath__GEN_15_0;
  assign _GEN_289 = dpath__GEN_289;
  assign _GEN_12_0 = cpath__GEN_12_1;
  assign _GEN_406 = cpath__GEN_406_0;
  assign _GEN_299 = dpath__GEN_299;
  assign _GEN_48 = cpath__GEN_48_0;
  assign _GEN_115 = cpath__GEN_115_0;
  assign _GEN_311 = dpath__GEN_311;
  assign _GEN_206 = dpath__GEN_206;
  assign _GEN_367 = dpath__GEN_367;
  assign _GEN_175 = dpath__GEN_175;
  assign _GEN_6_0 = cpath__GEN_6_1;
  assign _GEN_305 = dpath__GEN_305;
  assign _GEN_33 = cpath__GEN_33_0;
  assign _GEN_274 = dpath__GEN_274;
  assign _GEN_121 = cpath__GEN_121_0;
  assign _GEN_307 = cpath__GEN_307_0;
  assign _GEN_373 = dpath__GEN_373;
  assign _GEN_375 = cpath__GEN_375_0;
  assign _GEN_229 = cpath__GEN_229_0;
  assign _GEN_94 = cpath__GEN_94_0;
  assign _GEN_292 = cpath__GEN_292_0;
  assign _GEN_183 = cpath__GEN_183_0;
  assign _GEN_376 = dpath__GEN_376;
  assign _GEN_382 = dpath__GEN_382;
  assign _GEN_0_0 = cpath__GEN_0_1;
  assign _GEN_10 = frontend__GEN_10_0;
  assign _GEN_370 = dpath__GEN_370;
  assign _GEN_349 = dpath__GEN_349;
  assign _GEN_196 = cpath__GEN_196_0;
  assign _GEN_186 = cpath__GEN_186_0;
  assign _GEN_262 = dpath__GEN_262;
  assign _GEN_400 = cpath__GEN_400_0;
  assign _GEN_103 = cpath__GEN_103_0;
  assign _GEN_264 = cpath__GEN_264_0;
  assign _GEN_295 = cpath__GEN_295_0;
  assign _GEN_355 = dpath__GEN_355;
  assign _GEN_159 = cpath__GEN_159_0;
  assign _GEN_202 = cpath__GEN_202_0;
  assign _GEN_171 = cpath__GEN_171_0;
  assign _GEN_357 = cpath__GEN_357_0;
  assign _GEN_270 = cpath__GEN_270_0;
  assign _GEN_277 = dpath__GEN_277;
  assign _GEN_384 = cpath__GEN_384_0;
  assign _GEN_36 = cpath__GEN_36_0;
  assign _GEN_285 = cpath__GEN_285_0;
  assign _GEN_165 = cpath__GEN_165_0;
  assign _GEN_279 = cpath__GEN_279_0;
  assign _GEN_194 = dpath__GEN_194;
  assign _GEN_184 = dpath__GEN_184;
  assign _GEN_378 = cpath__GEN_378_0;
  assign _GEN_293 = dpath__GEN_293;
  assign _GEN_21_0 = cpath__GEN_21_1;
  assign _GEN_301 = cpath__GEN_301_0;
  assign _GEN_157 = dpath__GEN_157;
  assign _GEN_3_0 = dpath__GEN_3_1;
  assign _GEN_361 = dpath__GEN_361;
  assign _GEN_394 = cpath__GEN_394_0;
  assign _GEN_15_0 = cpath__GEN_15_1;
  assign _GEN_256 = dpath__GEN_256;
  assign _GEN_363 = cpath__GEN_363_0;
  assign _GEN_9_2 = cpath__GEN_9_3;
  assign _GEN_258 = cpath__GEN_258_0;
  assign _GEN_97 = cpath__GEN_97_0;
  assign _GEN_283 = dpath__GEN_283;
  assign _GEN_163 = dpath__GEN_163;
  assign _GEN_178 = dpath__GEN_178;
  assign _GEN_345 = cpath__GEN_345_0;
  assign _GEN_339 = cpath__GEN_339_0;
  assign _GEN_8 = dpath__GEN_8_0;
  assign _GEN_11 = dpath__GEN_11_0;
  assign _GEN_18 = cpath__GEN_18_0;
  assign _GEN_259 = dpath__GEN_259;
  assign _GEN_147 = cpath__GEN_147_0;
  assign _GEN_358 = dpath__GEN_358;
  assign _GEN_330 = cpath__GEN_330_0;
  assign _GEN_172 = dpath__GEN_172;
  assign _GEN_86 = cpath__GEN_86_0;
  assign _GEN_13 = frontend__GEN_13_0;
  assign _GEN_271 = dpath__GEN_271;
  assign _GEN_265 = dpath__GEN_265;
  assign _GEN_280 = dpath__GEN_280;
  assign _GEN_160 = dpath__GEN_160;
  assign _GEN_273 = cpath__GEN_273_0;
  assign _GEN_343 = dpath__GEN_343;
  assign _GEN_379 = dpath__GEN_379;
  assign _GEN_351 = cpath__GEN_351_0;
  assign _GEN_238 = dpath__GEN_238;
  assign _GEN_231 = cpath__GEN_231_0;
  assign _GEN_189 = cpath__GEN_189_0;
  assign _GEN_337 = dpath__GEN_337;
  assign _GEN_153 = cpath__GEN_153_0;
  assign _GEN_288 = cpath__GEN_288_0;
  assign _GEN_364 = dpath__GEN_364;
  assign _GEN_244 = dpath__GEN_244;
  assign _GEN_366 = cpath__GEN_366_0;
  assign _GEN_252 = cpath__GEN_252_0;
  assign _GEN_180 = cpath__GEN_180_0;
  assign _GEN_166 = dpath__GEN_166;
  assign _GEN_71 = cpath__GEN_71_0;
  assign _GEN_174 = cpath__GEN_174_0;
  assign _GEN_168 = cpath__GEN_168_0;
  assign _GEN_372 = cpath__GEN_372_0;
  assign _GEN_3_1 = cpath__GEN_3_2;
  assign _GEN_387 = cpath__GEN_387_0;
  assign _GEN_246 = cpath__GEN_246_0;
  assign _GEN_267 = cpath__GEN_267_0;
  assign _GEN_286 = dpath__GEN_286;
  assign _GEN_151 = dpath__GEN_151;
  assign _GEN_187 = dpath__GEN_187;
  assign _GEN_354 = cpath__GEN_354_0;
  assign _GEN_213 = cpath__GEN_213_0;
  assign _GEN_249 = cpath__GEN_249_0;
  assign _GEN_319_0 = dpath__GEN_319_0;
  assign _GEN_268 = dpath__GEN_268;
  assign _GEN_240 = cpath__GEN_240_0;
  assign _GEN_141 = cpath__GEN_141_0;
  assign _GEN_135 = cpath__GEN_135_0;
  assign _GEN_226_0 = dpath__GEN_226_0;
  assign _GEN_234 = cpath__GEN_234_0;
  assign _GEN_348 = cpath__GEN_348_0;
  assign _GEN_261 = cpath__GEN_261_0;
  assign _GEN_312 = cpath__GEN_312_0;
  assign _GEN_53 = cpath__GEN_53_0;
  assign _GEN_333 = cpath__GEN_333_0;
  assign _GEN_147_0 = dpath__GEN_147_0;
  assign _GEN_68 = cpath__GEN_68_0;
  assign _GEN_156 = cpath__GEN_156_0;
  assign _GEN_352 = dpath__GEN_352;
  assign _GEN_247_0 = dpath__GEN_247_0;
  assign _GEN_360 = cpath__GEN_360_0;
  assign _GEN_369 = cpath__GEN_369_0;
  assign _GEN_325_0 = dpath__GEN_325_0;
  assign _GEN_2 = dpath__GEN_2_0;
  assign _GEN_74 = cpath__GEN_74_0;
  assign _GEN_327 = cpath__GEN_327_0;
  assign _GEN_169 = dpath__GEN_169;
  assign _GEN_89 = cpath__GEN_89_0;
  assign _GEN_162 = cpath__GEN_162_0;
  assign _GEN_232_0 = dpath__GEN_232_0;
  assign _GEN_426 = cpath__GEN_426_0;
  assign _GEN_7_0 = frontend__GEN_7_1;
  assign _GEN_331_0 = dpath__GEN_331_0;
  assign _GEN_129 = cpath__GEN_129_0;
  assign _GEN_346 = dpath__GEN_346;
  assign _GEN_154 = dpath__GEN_154;
  assign _GEN_340 = dpath__GEN_340;
  assign _GEN_253 = dpath__GEN_253;
  assign _GEN_228 = cpath__GEN_228_0;
  assign _GEN_411 = cpath__GEN_411_0;
  assign _GEN_255 = cpath__GEN_255_0;
  assign _GEN_120 = cpath__GEN_120_0;
  assign _GEN_211_0 = dpath__GEN_211_0;
  assign _GEN_80 = cpath__GEN_80_0;
  assign _GEN_220_0 = dpath__GEN_220_0;
  assign _GEN_342 = cpath__GEN_342_0;
  assign _GEN_229_0 = dpath__GEN_229_0;
  assign _GEN_393 = cpath__GEN_393_0;
  assign _GEN_292_0 = dpath__GEN_292_0;
  assign _GEN_307_0 = dpath__GEN_307_0;
  assign _GEN_193_0 = dpath__GEN_193_0;
  assign _GEN_56 = cpath__GEN_56_0;
  assign _GEN_144 = cpath__GEN_144_0;
  assign _GEN_17 = dpath__GEN_17_0;
  assign _GEN_11_1 = dpath__GEN_11_2;
  assign _GEN_408 = cpath__GEN_408_0;
  assign _GEN_222 = cpath__GEN_222_0;
  assign _GEN_313_0 = dpath__GEN_313_0;
  assign _GEN_117 = cpath__GEN_117_0;
  assign _GEN_328 = dpath__GEN_328;
  assign _GEN_321 = cpath__GEN_321_0;
  assign _GEN_2_0 = dpath__GEN_2_1;
  assign _GEN_235 = dpath__GEN_235;
  assign _GEN_243 = cpath__GEN_243_0;
  assign _GEN_237 = cpath__GEN_237_0;
  assign _GEN_123 = cpath__GEN_123_0;
  assign _GEN_102 = cpath__GEN_102_0;
  assign _GEN_3_2 = dpath__GEN_3_3;
  assign _GEN_62 = cpath__GEN_62_0;
  assign _GEN_150 = cpath__GEN_150_0;
  assign _GEN_336 = cpath__GEN_336_0;
  assign _GEN_201 = cpath__GEN_201_0;
  assign _GEN_195 = cpath__GEN_195_0;
  assign _GEN_23 = dpath__GEN_23_0;
  assign _GEN_414 = cpath__GEN_414_0;
  assign _GEN_250 = dpath__GEN_250;
  assign _GEN_300 = cpath__GEN_300_0;
  assign _GEN_294 = cpath__GEN_294_0;
  assign _GEN_309 = cpath__GEN_309_0;
  assign _GEN_77 = cpath__GEN_77_0;
  assign _GEN_208_0 = dpath__GEN_208_0;
  assign _GEN_83 = cpath__GEN_83_0;
  assign _GEN_214_0 = dpath__GEN_214_0;
  assign _GEN_216 = cpath__GEN_216_0;
  assign _GEN_241 = dpath__GEN_241;
  assign _GEN_420 = cpath__GEN_420_0;
  assign _GEN_35 = cpath__GEN_35_0;
  assign _GEN_5_0 = dpath__GEN_5_1;
  assign _GEN_41 = cpath__GEN_41_0;
  assign _GEN_315 = cpath__GEN_315_0;
  assign _GEN_429 = cpath__GEN_429_0;
  assign _GEN_138 = cpath__GEN_138_0;
  assign _GEN_334 = dpath__GEN_334;
  assign _GEN_217 = dpath__GEN_217;
  assign _GEN_402 = cpath__GEN_402_0;
  assign _GEN_17_0 = cpath__GEN_17_1;
  assign _GEN_225 = cpath__GEN_225_0;
  assign _GEN_105 = cpath__GEN_105_0;
  assign _GEN_316 = dpath__GEN_316;
  assign _GEN_50 = cpath__GEN_50_0;
  assign _GEN_44 = cpath__GEN_44_0;
  assign _GEN_324 = cpath__GEN_324_0;
  assign _GEN_180_0 = dpath__GEN_180_0;
  assign _GEN_318 = cpath__GEN_318_0;
  assign _GEN_384_0 = dpath__GEN_384_0;
  assign _GEN_396 = cpath__GEN_396_0;
  assign _GEN_386 = cpath__GEN_386_0;
  assign _GEN_38 = cpath__GEN_38_0;
  assign _GEN_301_0 = dpath__GEN_301_0;
  assign _GEN_196_0 = dpath__GEN_196_0;
  assign _GEN_186_0 = dpath__GEN_186_0;
  assign _GEN_65 = cpath__GEN_65_0;
  assign _GEN_295_0 = dpath__GEN_295_0;
  assign _GEN_20 = dpath__GEN_20_0;
  assign _GEN_223 = dpath__GEN_223;
  assign _GEN_23_0 = cpath__GEN_23_1;
  assign _GEN_417 = cpath__GEN_417_0;
  assign _GEN_111 = cpath__GEN_111_0;
  assign _GEN_322 = dpath__GEN_322;
  assign _GEN_210 = cpath__GEN_210_0;
  assign _GEN_5_1 = dpath__GEN_5_2;
  assign _GEN_219 = cpath__GEN_219_0;
  assign _GEN_279_0 = dpath__GEN_279_0;
  assign _GEN_310_0 = dpath__GEN_310_0;
  assign _GEN_285_0 = dpath__GEN_285_0;
  assign _GEN_423 = cpath__GEN_423_0;
  assign _GEN_132 = cpath__GEN_132_0;
  assign _GEN_126 = cpath__GEN_126_0;
  assign _GEN_287 = cpath__GEN_287_0;
  assign _GEN_202_0 = dpath__GEN_202_0;
  assign _GEN_378_0 = dpath__GEN_378_0;
  assign _GEN_90 = cpath__GEN_90_0;
  assign _GEN_204 = cpath__GEN_204_0;
  assign _GEN_99 = cpath__GEN_99_0;
  assign _GEN_303 = cpath__GEN_303_0;
  assign _GEN_297 = cpath__GEN_297_0;
  assign _GEN_59 = cpath__GEN_59_0;
  assign _GEN_188 = cpath__GEN_188_0;
  assign _GEN_198 = cpath__GEN_198_0;
  assign _GEN_351_0 = dpath__GEN_351_0;
  assign _GEN_176 = cpath__GEN_176_0;
  assign _GEN_387_0 = dpath__GEN_387_0;
  assign _GEN_11_2 = cpath__GEN_11_3;
  assign _GEN_380 = cpath__GEN_380_0;
  assign _GEN_93 = cpath__GEN_93_0;
  assign _GEN_161 = cpath__GEN_161_0;
  assign _GEN_192 = cpath__GEN_192_0;
  assign _GEN_189_0 = dpath__GEN_189_0;
  assign _GEN_14_0 = dpath__GEN_14_1;
  assign _GEN_372_0 = dpath__GEN_372_0;
  assign _GEN_207 = cpath__GEN_207_0;
  assign _GEN_267_0 = dpath__GEN_267_0;
  assign _GEN_405 = cpath__GEN_405_0;
  assign _GEN_260 = cpath__GEN_260_0;
  assign _GEN_26 = cpath__GEN_26_0;
  assign _GEN_114 = cpath__GEN_114_0;
  assign _GEN_269 = cpath__GEN_269_0;
  assign _GEN_174_0 = dpath__GEN_174_0;
  assign _GEN_205_0 = dpath__GEN_205_0;
  assign _GEN_182 = cpath__GEN_182_0;
  assign _GEN_399 = cpath__GEN_399_0;
  assign _GEN_368 = cpath__GEN_368_0;
  assign _GEN_273_0 = dpath__GEN_273_0;
  assign _GEN_390 = cpath__GEN_390_0;
  assign _GEN_32 = cpath__GEN_32_0;
  assign _GEN_281 = cpath__GEN_281_0;
  assign _GEN_275 = cpath__GEN_275_0;
  assign _GEN_291 = cpath__GEN_291_0;
  assign _GEN_168_0 = dpath__GEN_168_0;
  assign _GEN_47 = cpath__GEN_47_0;
  assign _GEN_199_0 = dpath__GEN_199_0;
  assign _GEN_5_2 = cpath__GEN_5_3;
  assign _GEN_389 = cpath__GEN_389_0;
  assign _GEN_298_0 = dpath__GEN_298_0;
  assign _GEN_304_0 = dpath__GEN_304_0;
  assign _GEN_306 = cpath__GEN_306_0;
  assign _GEN_366_0 = dpath__GEN_366_0;
  assign _GEN_8_1 = dpath__GEN_8_2;
  assign _GEN_374 = cpath__GEN_374_0;
  assign _GEN_108 = cpath__GEN_108_0;
  assign _GEN_360_0 = dpath__GEN_360_0;
  assign _GEN_288_0 = dpath__GEN_288_0;
  assign _GEN_356 = cpath__GEN_356_0;
  assign _GEN_375_0 = dpath__GEN_375_0;
  assign _GEN_255_0 = dpath__GEN_255_0;
  assign _GEN_261_0 = dpath__GEN_261_0;
  assign _GEN_20_0 = cpath__GEN_20_1;
  assign _GEN_14_1 = cpath__GEN_14_2;
  assign _GEN_29 = cpath__GEN_29_0;
  assign _GEN_270_0 = dpath__GEN_270_0;
  assign _GEN_150_0 = dpath__GEN_150_0;
  assign _GEN_333_0 = dpath__GEN_333_0;
  assign _GEN_82 = cpath__GEN_82_0;
  assign _GEN_177_0 = dpath__GEN_177_0;
  assign _GEN_170 = cpath__GEN_170_0;
  assign _GEN_381_0 = dpath__GEN_381_0;
  assign _GEN_185 = cpath__GEN_185_0;
  assign _GEN_1_1 = dpath__GEN_1_2;
  assign _GEN_276_0 = dpath__GEN_276_0;
  assign _GEN_10_0 = dpath__GEN_10_1;
  assign _GEN_278 = cpath__GEN_278_0;
  assign _GEN_143 = cpath__GEN_143_0;
  assign _GEN_354_0 = dpath__GEN_354_0;
  assign _GEN_348_0 = dpath__GEN_348_0;
  assign _GEN_249_0 = dpath__GEN_249_0;
  assign _GEN_96 = cpath__GEN_96_0;
  assign _GEN_9_3 = frontend__GEN_9_4;
  assign _GEN_263 = cpath__GEN_263_0;
  assign _GEN_164 = cpath__GEN_164_0;
  assign _GEN_158 = cpath__GEN_158_0;
  assign _GEN_369_0 = dpath__GEN_369_0;
  assign _GEN_183_0 = dpath__GEN_183_0;
  assign _GEN_362 = cpath__GEN_362_0;
  assign _GEN_377 = cpath__GEN_377_0;
  assign _GEN_257 = cpath__GEN_257_0;
  assign _GEN_282_0 = dpath__GEN_282_0;
  assign _GEN_284 = cpath__GEN_284_0;
  assign _GEN_179 = cpath__GEN_179_0;
  assign _GEN_383 = cpath__GEN_383_0;
  assign _GEN_242 = cpath__GEN_242_0;
  assign _GEN_8_2 = cpath__GEN_8_3;
  assign _GEN_162_0 = dpath__GEN_162_0;
  assign _GEN_156_0 = dpath__GEN_156_0;
  assign _GEN_341 = cpath__GEN_341_0;
  assign _GEN_76 = cpath__GEN_76_0;
  assign _GEN_165_0 = dpath__GEN_165_0;
  assign _GEN_173 = cpath__GEN_173_0;
  assign _GEN_224_0 = cpath__GEN_224_1;
  assign _GEN_359 = cpath__GEN_359_0;
  assign _GEN_251 = cpath__GEN_251_0;
  assign _GEN_131 = cpath__GEN_131_0;
  assign _GEN_7_1 = dpath__GEN_7_2;
  assign _GEN_146 = cpath__GEN_146_0;
  assign _GEN_342_0 = dpath__GEN_342_0;
  assign _GEN_350 = cpath__GEN_350_0;
  assign _GEN_344 = cpath__GEN_344_0;
  assign _GEN_239_0 = cpath__GEN_239_1;
  assign _GEN_264_0 = dpath__GEN_264_0;
  assign _GEN_272 = cpath__GEN_272_0;
  assign _GEN_64 = cpath__GEN_64_0;
  assign _GEN_58 = cpath__GEN_58_0;
  assign _GEN_159_0 = dpath__GEN_159_0;
  assign _GEN_222_0 = dpath__GEN_222_0;
  assign _GEN_363_0 = dpath__GEN_363_0;
  assign _GEN_357_0 = dpath__GEN_357_0;
  assign _GEN_230 = cpath__GEN_230_0;
  assign _GEN_365 = cpath__GEN_365_0;
  assign _GEN_321_0 = dpath__GEN_321_0;
  assign _GEN_7_2 = dpath__GEN_7_3;
  assign _GEN_330_0 = dpath__GEN_330_0;
  assign _GEN_323_0 = cpath__GEN_323_1;
  assign _GEN_85 = cpath__GEN_85_0;
  assign _GEN_338_0 = cpath__GEN_338_1;
  assign _GEN_79 = cpath__GEN_79_0;
  assign _GEN_243_0 = dpath__GEN_243_0;
  assign _GEN_2_2 = cpath__GEN_2_3;
  assign _GEN_237_0 = dpath__GEN_237_0;
  assign _GEN_245 = cpath__GEN_245_0;
  assign _GEN_12_1 = frontend__GEN_12_2;
  assign _GEN_315_0 = dpath__GEN_315_0;
  assign _GEN_336_0 = dpath__GEN_336_0;
  assign _GEN_70 = cpath__GEN_70_0;
  assign _GEN_152 = cpath__GEN_152_0;
  assign _GEN_167 = cpath__GEN_167_0;
  assign _GEN_422 = cpath__GEN_422_0;
  assign _GEN_258_0 = dpath__GEN_258_0;
  assign _GEN_371 = cpath__GEN_371_0;
  assign _GEN_266 = cpath__GEN_266_0;
  assign _GEN_125 = cpath__GEN_125_0;
  assign _GEN_171_0 = dpath__GEN_171_0;
  assign _GEN_212_0 = cpath__GEN_212_1;
  assign _GEN_303_0 = dpath__GEN_303_0;
  assign _GEN_254 = cpath__GEN_254_0;
  assign _GEN_146_0 = dpath__GEN_146_0;
  assign _GEN_13_0 = dpath__GEN_13_1;
  assign _GEN_155 = cpath__GEN_155_0;
  assign _GEN_149 = cpath__GEN_149_0;
  assign _GEN_225_0 = dpath__GEN_225_0;
  assign _GEN_227 = cpath__GEN_227_0;
  assign _GEN_113 = cpath__GEN_113_0;
  assign _GEN_140 = cpath__GEN_140_0;
  assign _GEN_326 = cpath__GEN_326_0;
  assign _GEN_7_3 = dpath__GEN_7_4;
  assign _GEN_231_0 = dpath__GEN_231_0;
  assign _GEN_425 = cpath__GEN_425_0;
  assign _GEN_404 = cpath__GEN_404_0;
  assign _GEN_240_0 = dpath__GEN_240_0;
  assign _GEN_353 = cpath__GEN_353_0;
  assign _GEN_248 = cpath__GEN_248_0;
  assign _GEN_107 = cpath__GEN_107_0;
  assign _GEN_6_3 = frontend__GEN_6_4;
  assign _GEN_311_0 = cpath__GEN_311_1;
  assign _GEN_339_0 = dpath__GEN_339_0;
  assign _GEN_153_0 = dpath__GEN_153_0;
  assign _GEN_73 = cpath__GEN_73_0;
  assign _GEN_67 = cpath__GEN_67_0;
  assign _GEN_347 = cpath__GEN_347_0;
  assign _GEN_206_0 = cpath__GEN_206_1;
  assign _GEN_252_0 = dpath__GEN_252_0;
  assign _GEN_410 = cpath__GEN_410_0;
  assign _GEN_297_0 = dpath__GEN_297_0;
  assign _GEN_419 = cpath__GEN_419_0;
  assign _GEN_233 = cpath__GEN_233_0;
  assign _GEN_305_0 = cpath__GEN_305_1;
  assign _GEN_128 = cpath__GEN_128_0;
  assign _GEN_324_0 = dpath__GEN_324_0;
  assign _GEN_332 = cpath__GEN_332_0;
  assign _GEN_219_0 = dpath__GEN_219_0;
  assign _GEN_88 = cpath__GEN_88_0;
  assign _GEN_1_3 = dpath__GEN_1_4;
  assign _GEN_246_0 = dpath__GEN_246_0;
  assign _GEN_318_0 = dpath__GEN_318_0;
  assign _GEN_52 = cpath__GEN_52_0;
  assign _GEN_46 = cpath__GEN_46_0;
  assign _GEN_134 = cpath__GEN_134_0;
  assign _GEN_345_0 = dpath__GEN_345_0;
  assign _GEN_204_0 = dpath__GEN_204_0;
  assign _GEN_213_0 = dpath__GEN_213_0;
  assign _GEN_228_0 = dpath__GEN_228_0;
  assign _GEN_221 = cpath__GEN_221_0;
  assign _GEN_407 = cpath__GEN_407_0;
  assign _GEN_382_0 = cpath__GEN_382_1;
  assign _GEN_28 = cpath__GEN_28_0;
  assign _GEN_281_0 = dpath__GEN_281_0;
  assign _GEN_4_1 = dpath__GEN_4_2;
  assign _GEN_40 = cpath__GEN_40_0;
  assign _GEN_55 = cpath__GEN_55_0;
  assign _GEN_329 = cpath__GEN_329_0;
  assign _GEN_194_0 = cpath__GEN_194_1;
  assign _GEN_392 = cpath__GEN_392_0;
  assign _GEN_0_2 = dpath__GEN_0_3;
  assign _GEN_234_0 = dpath__GEN_234_0;
  assign _GEN_10_2 = dpath__GEN_10_3;
  assign _GEN_236 = cpath__GEN_236_0;
  assign _GEN_101 = cpath__GEN_101_0;
  assign _GEN_312_0 = dpath__GEN_312_0;
  assign _GEN_192_0 = dpath__GEN_192_0;
  assign _GEN_306_0 = dpath__GEN_306_0;
  assign _GEN_61 = cpath__GEN_61_0;
  assign _GEN_207_0 = dpath__GEN_207_0;
  assign _GEN_16 = dpath__GEN_16_0;
  assign _GEN_22 = dpath__GEN_22_0;
  assign _GEN_300_0 = dpath__GEN_300_0;
  assign _GEN_34 = cpath__GEN_34_0;
  assign _GEN_116 = cpath__GEN_116_0;
  assign _GEN_122 = cpath__GEN_122_0;
  assign _GEN_327_0 = dpath__GEN_327_0;
  assign _GEN_182_0 = dpath__GEN_182_0;
  assign _GEN_320_0 = cpath__GEN_320_1;
  assign _GEN_215 = cpath__GEN_215_0;
  assign _GEN_335 = cpath__GEN_335_0;
  assign _GEN_291_0 = dpath__GEN_291_0;
  assign _GEN_290 = dpath__GEN_290;
  assign _GEN_293_0 = cpath__GEN_293_1;
  assign _GEN_428 = cpath__GEN_428_0;
  assign _GEN_49 = cpath__GEN_49_0;
  assign _GEN_137 = cpath__GEN_137_0;
  assign _GEN_200_0 = cpath__GEN_200_1;
  assign _GEN_209 = cpath__GEN_209_0;
  assign _GEN_95 = cpath__GEN_95_0;
  assign _GEN_413 = cpath__GEN_413_0;
  assign _GEN_314 = cpath__GEN_314_0;
  assign _GEN_308 = cpath__GEN_308_0;
  assign _GEN_4_2 = dpath__GEN_4_3;
  assign _GEN_383_0 = dpath__GEN_383_0;
  assign _GEN_16_0 = cpath__GEN_16_1;
  assign _GEN_395 = cpath__GEN_395_0;
  assign _GEN_385_0 = cpath__GEN_385_1;
  assign _GEN_104 = cpath__GEN_104_0;
  assign _GEN_195_0 = dpath__GEN_195_0;
  assign _GEN_302_0 = cpath__GEN_302_1;
  assign _GEN_317_0 = cpath__GEN_317_1;
  assign _GEN_203_0 = cpath__GEN_203_1;
  assign _GEN_172_0 = cpath__GEN_172_1;
  assign _GEN_197_0 = cpath__GEN_197_1;
  assign _GEN_370_0 = cpath__GEN_370_1;
  assign _GEN_416 = cpath__GEN_416_0;
  assign _GEN_22_0 = cpath__GEN_22_1;
  assign _GEN_271_0 = cpath__GEN_271_1;
  assign _GEN_119 = cpath__GEN_119_0;
  assign _GEN_185_0 = dpath__GEN_185_0;
  assign _GEN_179_0 = dpath__GEN_179_0;
  assign _GEN_216_0 = dpath__GEN_216_0;
  assign _GEN_379_0 = cpath__GEN_379_1;
  assign _GEN_187_0 = cpath__GEN_187_1;
  assign _GEN_401 = cpath__GEN_401_0;
  assign _GEN_43 = cpath__GEN_43_0;
  assign _GEN_278_0 = dpath__GEN_278_0;
  assign _GEN_296_0 = cpath__GEN_296_1;
  assign _GEN_286_0 = cpath__GEN_286_1;
  assign _GEN_201_0 = dpath__GEN_201_0;
  assign _GEN_364_0 = cpath__GEN_364_1;
  assign _GEN_1_4 = cpath__GEN_1_5;
  assign _GEN_210_0 = dpath__GEN_210_0;
  assign _GEN_98 = cpath__GEN_98_0;
  assign _GEN_263_0 = dpath__GEN_263_0;
  assign _GEN_309_0 = dpath__GEN_309_0;
  assign _GEN_37 = cpath__GEN_37_0;
  assign _GEN_164_0 = dpath__GEN_164_0;
  assign _GEN_110 = cpath__GEN_110_0;
  assign _GEN_362_0 = dpath__GEN_362_0;
  assign _GEN_19 = dpath__GEN_19_0;
  assign _GEN_377_0 = dpath__GEN_377_0;
  assign _GEN_218_0 = cpath__GEN_218_1;
  assign _GEN_294_0 = dpath__GEN_294_0;
  assign _GEN_284_0 = dpath__GEN_284_0;
  assign _GEN_371_0 = dpath__GEN_371_0;
  assign _GEN_260_0 = dpath__GEN_260_0;
  assign _GEN_266_0 = dpath__GEN_266_0;
  assign _GEN_380_0 = dpath__GEN_380_0;
  assign _GEN_25 = cpath__GEN_25_0;
  assign _GEN_365_0 = dpath__GEN_365_0;
  assign _GEN_181_0 = cpath__GEN_181_1;
  assign _GEN_175_0 = cpath__GEN_175_1;
  assign _GEN_251_0 = dpath__GEN_251_0;
  assign _GEN_15_1 = dpath__GEN_15_2;
  assign _GEN_289_0 = cpath__GEN_289_1;
  assign _GEN_359_0 = dpath__GEN_359_0;
  assign _GEN_352_0 = cpath__GEN_352_1;
  assign _GEN_14_2 = frontend__GEN_14_3;
  assign _GEN_152_0 = dpath__GEN_152_0;
  assign _GEN_31 = cpath__GEN_31_0;
  assign _GEN_274_0 = cpath__GEN_274_1;
  assign _GEN_160_0 = cpath__GEN_160_1;
  assign _GEN_169_0 = cpath__GEN_169_1;
  assign _GEN_191_0 = cpath__GEN_191_1;
  assign _GEN_188_0 = dpath__GEN_188_0;
  assign _GEN_373_0 = cpath__GEN_373_1;
  assign _GEN_19_0 = cpath__GEN_19_1;
  assign _GEN_367_0 = cpath__GEN_367_1;
  assign _GEN_268_0 = cpath__GEN_268_1;
  assign _GEN_173_0 = dpath__GEN_173_0;
  assign _GEN_290_0 = cpath__GEN_290_1;
  assign _GEN_280_0 = cpath__GEN_280_1;
  assign _GEN_287_0 = dpath__GEN_287_0;
  assign _GEN_154_0 = cpath__GEN_154_1;
  assign _GEN_87 = cpath__GEN_87_0;
  assign _GEN_299_0 = cpath__GEN_299_1;
  assign _GEN_386_0 = dpath__GEN_386_0;
  assign _GEN_10_3 = cpath__GEN_10_4;
  assign _GEN_245_0 = dpath__GEN_245_0;
  assign _GEN_398 = cpath__GEN_398_0;
  assign _GEN_4_3 = cpath__GEN_4_4;
  assign _GEN_388_0 = cpath__GEN_388_1;
  assign _GEN_253_0 = cpath__GEN_253_1;
  assign _GEN_92 = cpath__GEN_92_0;
  assign _GEN_5_3 = frontend__GEN_5_4;
  assign _GEN_272_0 = dpath__GEN_272_0;
  assign _GEN_344_0 = dpath__GEN_344_0;
  assign _GEN_198_0 = dpath__GEN_198_0;
  assign _GEN_167_0 = dpath__GEN_167_0;
  assign _GEN_346_0 = cpath__GEN_346_1;
  assign _GEN_334_0 = cpath__GEN_334_1;
  assign _GEN_340_0 = cpath__GEN_340_1;
  assign _GEN_254_0 = dpath__GEN_254_0;
  assign _GEN_13_2 = cpath__GEN_13_3;
  assign _GEN_3_4 = dpath__GEN_3_5;
  assign _GEN_256_0 = cpath__GEN_256_1;
  assign _GEN_328_0 = cpath__GEN_328_1;
  assign _GEN_161_0 = dpath__GEN_161_0;
  assign _GEN_347_0 = dpath__GEN_347_0;
  assign _GEN_81 = cpath__GEN_81_0;
  assign _GEN_355_0 = cpath__GEN_355_1;
  assign _GEN_170_0 = dpath__GEN_170_0;
  assign _GEN_7_5 = cpath__GEN_7_6;
  assign _GEN_8_3 = frontend__GEN_8_4;
  assign _GEN_275_0 = dpath__GEN_275_0;
  assign _GEN_269_0 = dpath__GEN_269_0;
  assign _GEN_155_0 = dpath__GEN_155_0;
  assign _GEN_277_0 = cpath__GEN_277_1;
  assign _GEN_69 = cpath__GEN_69_0;
  assign _GEN_157_0 = cpath__GEN_157_1;
  assign _GEN_368_0 = dpath__GEN_368_0;
  assign _GEN_233_0 = dpath__GEN_233_0;
  assign _GEN_227_0 = dpath__GEN_227_0;
  assign _GEN_235_0 = cpath__GEN_235_1;
  assign _GEN_184_0 = cpath__GEN_184_1;
  assign _GEN_326_0 = dpath__GEN_326_0;
  assign _GEN_149_0 = dpath__GEN_149_0;
  assign _GEN_60 = cpath__GEN_60_0;
  assign _GEN_283_0 = cpath__GEN_283_1;
  assign _GEN_142 = cpath__GEN_142_0;
  assign _GEN_353_0 = dpath__GEN_353_0;
  assign _GEN_178_0 = cpath__GEN_178_1;
  assign _GEN_248_0 = dpath__GEN_248_0;
  assign _GEN_241_0 = cpath__GEN_241_1;
  assign _GEN_361_0 = cpath__GEN_361_1;
  assign _GEN_136 = cpath__GEN_136_0;
  assign _GEN_75 = cpath__GEN_75_0;
  assign _GEN_163_0 = cpath__GEN_163_1;
  assign _GEN_349_0 = cpath__GEN_349_1;
  assign _GEN_374_0 = dpath__GEN_374_0;
  assign _GEN_427 = cpath__GEN_427_0;
  assign _GEN_376_0 = cpath__GEN_376_1;
  assign _GEN_262_0 = cpath__GEN_262_1;
  assign _GEN_332_0 = dpath__GEN_332_0;
  assign _GEN_176_0 = dpath__GEN_176_0;
  assign _GEN_166_0 = cpath__GEN_166_1;
  assign _GEN_358_0 = cpath__GEN_358_1;
  assign _GEN_314_0 = dpath__GEN_314_0;
  assign _GEN_308_0 = dpath__GEN_308_0;
  assign _GEN_42 = cpath__GEN_42_0;
  assign _GEN_265_0 = cpath__GEN_265_1;
  assign _GEN_316_0 = cpath__GEN_316_1;
  assign _GEN_130 = cpath__GEN_130_0;
  assign _GEN_124 = cpath__GEN_124_0;
  assign _GEN_341_0 = dpath__GEN_341_0;
  assign _GEN_343_0 = cpath__GEN_343_1;
  assign _GEN_223_0 = cpath__GEN_223_1;
  assign _GEN_238_0 = cpath__GEN_238_1;
  assign _GEN_118 = cpath__GEN_118_0;
  assign _GEN_5_4 = dpath__GEN_5_5;
  assign _GEN_151_0 = cpath__GEN_151_1;
  assign _GEN_145 = cpath__GEN_145_0;
  assign _GEN_337_0 = cpath__GEN_337_1;
  assign _GEN_18_0 = dpath__GEN_18_1;
  assign _GEN_356_0 = dpath__GEN_356_0;
  assign _GEN_244_0 = cpath__GEN_244_1;
  assign _GEN_409 = cpath__GEN_409_0;
  assign _GEN_11_3 = frontend__GEN_11_4;
  assign _GEN_322_0 = cpath__GEN_322_1;
  assign _GEN_158_0 = dpath__GEN_158_0;
  assign _GEN_209_0 = dpath__GEN_209_0;
  assign _GEN_78 = cpath__GEN_78_0;
  assign _GEN_217_0 = cpath__GEN_217_1;
  assign _GEN_221_0 = dpath__GEN_221_0;
  assign _GEN_236_0 = dpath__GEN_236_0;
  assign _GEN_421 = cpath__GEN_421_0;
  assign _GEN_415 = cpath__GEN_415_0;
  assign _GEN_335_0 = dpath__GEN_335_0;
  assign _GEN_329_0 = dpath__GEN_329_0;
  assign _GEN_63 = cpath__GEN_63_0;
  assign _GEN_230_0 = dpath__GEN_230_0;
  assign _GEN_242_0 = dpath__GEN_242_0;
  assign _GEN_257_0 = dpath__GEN_257_0;
  assign _GEN_6_4 = dpath__GEN_6_5;
  assign _GEN_57 = cpath__GEN_57_0;
  assign _GEN_250_0 = cpath__GEN_250_1;
  assign _GEN_259_0 = cpath__GEN_259_1;
  assign _GEN_139 = cpath__GEN_139_0;
  assign _GEN_350_0 = dpath__GEN_350_0;
  assign _GEN_215_0 = dpath__GEN_215_0;
  assign _GEN_84 = cpath__GEN_84_0;
  assign frontend_clock = clock;
  assign frontend_reset = reset;
  assign frontend_io_cpu_req_valid = cpath_io_imem_req_valid;
  assign frontend_io_cpu_req_bits_pc = dpath_io_imem_req_bits_pc;
  assign frontend_io_cpu_resp_ready = dpath_io_imem_resp_ready;
  assign frontend_io_imem_resp_bits_data = io_imem_resp_bits_data;
  assign cpath_clock = clock;
  assign cpath_io_imem_resp_valid = frontend_io_cpu_resp_valid;
  assign cpath_io_imem_resp_bits_inst = frontend_io_cpu_resp_bits_inst;
  assign cpath_io_dat_br_eq = dpath_io_dat_br_eq;
  assign cpath_io_dat_br_lt = dpath_io_dat_br_lt;
  assign cpath_io_dat_br_ltu = dpath_io_dat_br_ltu;
  assign cpath_io_dat_csr_eret = dpath_io_dat_csr_eret;
  assign dpath_clock = clock;
  assign dpath_reset = reset;
  assign dpath_io_imem_resp_valid = frontend_io_cpu_resp_valid;
  assign dpath_io_imem_resp_bits_pc = frontend_io_cpu_resp_bits_pc;
  assign dpath_io_imem_resp_bits_inst = frontend_io_cpu_resp_bits_inst;
  assign dpath_io_dmem_resp_bits_data = io_dmem_resp_bits_data;
  assign dpath_io_ctl_exe_kill = cpath_io_ctl_exe_kill;
  assign dpath_io_ctl_pc_sel = cpath_io_ctl_pc_sel;
  assign dpath_io_ctl_brjmp_sel = cpath_io_ctl_brjmp_sel;
  assign dpath_io_ctl_op1_sel = cpath_io_ctl_op1_sel;
  assign dpath_io_ctl_op2_sel = cpath_io_ctl_op2_sel;
  assign dpath_io_ctl_alu_fun = cpath_io_ctl_alu_fun;
  assign dpath_io_ctl_wb_sel = cpath_io_ctl_wb_sel;
  assign dpath_io_ctl_rf_wen = cpath_io_ctl_rf_wen;
  assign dpath_io_ctl_bypassable = cpath_io_ctl_bypassable;
  assign dpath_io_ctl_csr_cmd = cpath_io_ctl_csr_cmd;
  assign dpath_io_ctl_dmem_fcn = cpath_io_ctl_dmem_fcn;
  assign dpath_io_ctl_dmem_typ = cpath_io_ctl_dmem_typ;
  assign dpath_io_ctl_exception = cpath_io_ctl_exception;
endmodule
module SyncMem( // @[:Sodor3Stage.fir@3768.2]
  input         metaReset,
  input         clock, // @[:Sodor3Stage.fir@3769.4]
  input  [20:0] io_dataInstr_0_addr, // @[:Sodor3Stage.fir@3771.4]
  output [31:0] io_dataInstr_0_data, // @[:Sodor3Stage.fir@3771.4]
  input  [20:0] io_dw_addr, // @[:Sodor3Stage.fir@3771.4]
  input  [31:0] io_dw_data, // @[:Sodor3Stage.fir@3771.4]
  input         io_dw_en, // @[:Sodor3Stage.fir@3771.4]
  output        _GEN_3_0,
  output        _GEN_2_2,
  output        _GEN_1_3,
  output        _GEN_0_4
);
  wire  mem_sparse_metaReset; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire  mem_sparse_clock; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire [20:0] mem_sparse_io_w_1_addr; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire  mem_sparse_io_w_1_en; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire [7:0] mem_sparse_io_w_1_data; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire [20:0] mem_sparse_io_r_0_addr; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire [7:0] mem_sparse_io_r_0_data; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire  mem_sparse_0_metaReset; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire  mem_sparse_0_clock; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire [20:0] mem_sparse_0_io_w_1_addr; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire  mem_sparse_0_io_w_1_en; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire [7:0] mem_sparse_0_io_w_1_data; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire [20:0] mem_sparse_0_io_r_0_addr; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire [7:0] mem_sparse_0_io_r_0_data; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire  mem_sparse_1_metaReset; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire  mem_sparse_1_clock; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire [20:0] mem_sparse_1_io_w_1_addr; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire  mem_sparse_1_io_w_1_en; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire [7:0] mem_sparse_1_io_w_1_data; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire [20:0] mem_sparse_1_io_r_0_addr; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire [7:0] mem_sparse_1_io_r_0_data; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire  mem_sparse_2_metaReset; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire  mem_sparse_2_clock; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire [20:0] mem_sparse_2_io_w_1_addr; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire  mem_sparse_2_io_w_1_en; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire [7:0] mem_sparse_2_io_w_1_data; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire [20:0] mem_sparse_2_io_r_0_addr; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire [7:0] mem_sparse_2_io_r_0_data; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  reg [20:0] underlying_0__T_54_addr_pipe_0;
  reg [31:0] _RAND_0;
  reg [20:0] underlying_1__T_54_addr_pipe_0;
  reg [31:0] _RAND_1;
  reg [20:0] underlying_2__T_54_addr_pipe_0;
  reg [31:0] _RAND_2;
  reg [20:0] underlying_3__T_54_addr_pipe_0;
  reg [31:0] _RAND_3;
  wire [7:0] underlying_1__T_54_data; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire [7:0] underlying_0__T_54_data; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire [15:0] _T_68; // @[memory.scala 82:55:Sodor3Stage.fir@3776.4]
  wire [7:0] underlying_3__T_54_data; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire [7:0] underlying_2__T_54_data; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  wire [15:0] _T_69; // @[memory.scala 82:55:Sodor3Stage.fir@3777.4]
  SparseMem_0 mem_sparse ( // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
    .metaReset(mem_sparse_metaReset),
    .clock(mem_sparse_clock),
    .io_w_1_addr(mem_sparse_io_w_1_addr),
    .io_w_1_en(mem_sparse_io_w_1_en),
    .io_w_1_data(mem_sparse_io_w_1_data),
    .io_r_0_addr(mem_sparse_io_r_0_addr),
    .io_r_0_data(mem_sparse_io_r_0_data)
  );
  SparseMem_0 mem_sparse_0 ( // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
    .metaReset(mem_sparse_0_metaReset),
    .clock(mem_sparse_0_clock),
    .io_w_1_addr(mem_sparse_0_io_w_1_addr),
    .io_w_1_en(mem_sparse_0_io_w_1_en),
    .io_w_1_data(mem_sparse_0_io_w_1_data),
    .io_r_0_addr(mem_sparse_0_io_r_0_addr),
    .io_r_0_data(mem_sparse_0_io_r_0_data)
  );
  SparseMem_0 mem_sparse_1 ( // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
    .metaReset(mem_sparse_1_metaReset),
    .clock(mem_sparse_1_clock),
    .io_w_1_addr(mem_sparse_1_io_w_1_addr),
    .io_w_1_en(mem_sparse_1_io_w_1_en),
    .io_w_1_data(mem_sparse_1_io_w_1_data),
    .io_r_0_addr(mem_sparse_1_io_r_0_addr),
    .io_r_0_data(mem_sparse_1_io_r_0_data)
  );
  SparseMem_0 mem_sparse_2 ( // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
    .metaReset(mem_sparse_2_metaReset),
    .clock(mem_sparse_2_clock),
    .io_w_1_addr(mem_sparse_2_io_w_1_addr),
    .io_w_1_en(mem_sparse_2_io_w_1_en),
    .io_w_1_data(mem_sparse_2_io_w_1_data),
    .io_r_0_addr(mem_sparse_2_io_r_0_addr),
    .io_r_0_data(mem_sparse_2_io_r_0_data)
  );
  assign mem_sparse_metaReset = metaReset;
  assign mem_sparse_0_metaReset = metaReset;
  assign mem_sparse_1_metaReset = metaReset;
  assign mem_sparse_2_metaReset = metaReset;
  assign underlying_1__T_54_data = mem_sparse_0_io_r_0_data; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  assign underlying_0__T_54_data = mem_sparse_io_r_0_data; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  assign _T_68 = {underlying_1__T_54_data,underlying_0__T_54_data}; // @[memory.scala 82:55:Sodor3Stage.fir@3776.4]
  assign underlying_3__T_54_data = mem_sparse_2_io_r_0_data; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  assign underlying_2__T_54_data = mem_sparse_1_io_r_0_data; // @[memory.scala 97:36:Sodor3Stage.fir@3773.4]
  assign _T_69 = {underlying_3__T_54_data,underlying_2__T_54_data}; // @[memory.scala 82:55:Sodor3Stage.fir@3777.4]
  assign io_dataInstr_0_data = {_T_69,_T_68};
  assign _GEN_3_0 = io_dw_en;
  assign _GEN_2_2 = io_dw_en;
  assign _GEN_1_3 = io_dw_en;
  assign _GEN_0_4 = io_dw_en;
  assign mem_sparse_clock = clock;
  assign mem_sparse_io_w_1_addr = io_dw_addr;
  assign mem_sparse_io_w_1_en = io_dw_en;
  assign mem_sparse_io_w_1_data = io_dw_data[7:0];
  assign mem_sparse_io_r_0_addr = underlying_0__T_54_addr_pipe_0;
  assign mem_sparse_0_clock = clock;
  assign mem_sparse_0_io_w_1_addr = io_dw_addr;
  assign mem_sparse_0_io_w_1_en = io_dw_en;
  assign mem_sparse_0_io_w_1_data = io_dw_data[15:8];
  assign mem_sparse_0_io_r_0_addr = underlying_1__T_54_addr_pipe_0;
  assign mem_sparse_1_clock = clock;
  assign mem_sparse_1_io_w_1_addr = io_dw_addr;
  assign mem_sparse_1_io_w_1_en = io_dw_en;
  assign mem_sparse_1_io_w_1_data = io_dw_data[23:16];
  assign mem_sparse_1_io_r_0_addr = underlying_2__T_54_addr_pipe_0;
  assign mem_sparse_2_clock = clock;
  assign mem_sparse_2_io_w_1_addr = io_dw_addr;
  assign mem_sparse_2_io_w_1_en = io_dw_en;
  assign mem_sparse_2_io_w_1_data = io_dw_data[31:24];
  assign mem_sparse_2_io_r_0_addr = underlying_3__T_54_addr_pipe_0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  underlying_0__T_54_addr_pipe_0 = _RAND_0[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  underlying_1__T_54_addr_pipe_0 = _RAND_1[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  underlying_2__T_54_addr_pipe_0 = _RAND_2[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  underlying_3__T_54_addr_pipe_0 = _RAND_3[20:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (metaReset) begin
      underlying_0__T_54_addr_pipe_0 <= 21'h0;
    end else begin
      underlying_0__T_54_addr_pipe_0 <= io_dataInstr_0_addr;
    end
    if (metaReset) begin
      underlying_1__T_54_addr_pipe_0 <= 21'h0;
    end else begin
      underlying_1__T_54_addr_pipe_0 <= io_dataInstr_0_addr;
    end
    if (metaReset) begin
      underlying_2__T_54_addr_pipe_0 <= 21'h0;
    end else begin
      underlying_2__T_54_addr_pipe_0 <= io_dataInstr_0_addr;
    end
    if (metaReset) begin
      underlying_3__T_54_addr_pipe_0 <= 21'h0;
    end else begin
      underlying_3__T_54_addr_pipe_0 <= io_dataInstr_0_addr;
    end
  end
endmodule
module SparseMem_0(
  input         metaReset,
  input         clock,
  input  [20:0] io_w_1_addr,
  input         io_w_1_en,
  input  [7:0]  io_w_1_data,
  input  [20:0] io_r_0_addr,
  output [7:0]  io_r_0_data
);
  reg [7:0] mem [0:31];
  reg [31:0] _RAND_0;
  wire [7:0] mem__T_959_data;
  wire [4:0] mem__T_959_addr;
  wire [7:0] mem__T_1124_data;
  wire [4:0] mem__T_1124_addr;
  wire [7:0] mem__T_1289_data;
  wire [4:0] mem__T_1289_addr;
  wire [7:0] mem__T_1484_data;
  wire [4:0] mem__T_1484_addr;
  wire  mem__T_1484_mask;
  wire  mem__T_1484_en;
  wire [7:0] mem__T_1670_data;
  wire [4:0] mem__T_1670_addr;
  wire  mem__T_1670_mask;
  wire  mem__T_1670_en;
  wire [4:0] _GEN_395;
  wire [4:0] _GEN_404;
  reg  addresses_0_valid;
  reg [31:0] _RAND_1;
  reg [20:0] addresses_0_bits;
  reg [31:0] _RAND_2;
  reg  addresses_1_valid;
  reg [31:0] _RAND_3;
  reg [20:0] addresses_1_bits;
  reg [31:0] _RAND_4;
  reg  addresses_2_valid;
  reg [31:0] _RAND_5;
  reg [20:0] addresses_2_bits;
  reg [31:0] _RAND_6;
  reg  addresses_3_valid;
  reg [31:0] _RAND_7;
  reg [20:0] addresses_3_bits;
  reg [31:0] _RAND_8;
  reg  addresses_4_valid;
  reg [31:0] _RAND_9;
  reg [20:0] addresses_4_bits;
  reg [31:0] _RAND_10;
  reg  addresses_5_valid;
  reg [31:0] _RAND_11;
  reg [20:0] addresses_5_bits;
  reg [31:0] _RAND_12;
  reg  addresses_6_valid;
  reg [31:0] _RAND_13;
  reg [20:0] addresses_6_bits;
  reg [31:0] _RAND_14;
  reg  addresses_7_valid;
  reg [31:0] _RAND_15;
  reg [20:0] addresses_7_bits;
  reg [31:0] _RAND_16;
  reg  addresses_8_valid;
  reg [31:0] _RAND_17;
  reg [20:0] addresses_8_bits;
  reg [31:0] _RAND_18;
  reg  addresses_9_valid;
  reg [31:0] _RAND_19;
  reg [20:0] addresses_9_bits;
  reg [31:0] _RAND_20;
  reg  addresses_10_valid;
  reg [31:0] _RAND_21;
  reg [20:0] addresses_10_bits;
  reg [31:0] _RAND_22;
  reg  addresses_11_valid;
  reg [31:0] _RAND_23;
  reg [20:0] addresses_11_bits;
  reg [31:0] _RAND_24;
  reg  addresses_12_valid;
  reg [31:0] _RAND_25;
  reg [20:0] addresses_12_bits;
  reg [31:0] _RAND_26;
  reg  addresses_13_valid;
  reg [31:0] _RAND_27;
  reg [20:0] addresses_13_bits;
  reg [31:0] _RAND_28;
  reg  addresses_14_valid;
  reg [31:0] _RAND_29;
  reg [20:0] addresses_14_bits;
  reg [31:0] _RAND_30;
  reg  addresses_15_valid;
  reg [31:0] _RAND_31;
  reg [20:0] addresses_15_bits;
  reg [31:0] _RAND_32;
  reg  addresses_16_valid;
  reg [31:0] _RAND_33;
  reg [20:0] addresses_16_bits;
  reg [31:0] _RAND_34;
  reg  addresses_17_valid;
  reg [31:0] _RAND_35;
  reg [20:0] addresses_17_bits;
  reg [31:0] _RAND_36;
  reg  addresses_18_valid;
  reg [31:0] _RAND_37;
  reg [20:0] addresses_18_bits;
  reg [31:0] _RAND_38;
  reg  addresses_19_valid;
  reg [31:0] _RAND_39;
  reg [20:0] addresses_19_bits;
  reg [31:0] _RAND_40;
  reg  addresses_20_valid;
  reg [31:0] _RAND_41;
  reg [20:0] addresses_20_bits;
  reg [31:0] _RAND_42;
  reg  addresses_21_valid;
  reg [31:0] _RAND_43;
  reg [20:0] addresses_21_bits;
  reg [31:0] _RAND_44;
  reg  addresses_22_valid;
  reg [31:0] _RAND_45;
  reg [20:0] addresses_22_bits;
  reg [31:0] _RAND_46;
  reg  addresses_23_valid;
  reg [31:0] _RAND_47;
  reg [20:0] addresses_23_bits;
  reg [31:0] _RAND_48;
  reg  addresses_24_valid;
  reg [31:0] _RAND_49;
  reg [20:0] addresses_24_bits;
  reg [31:0] _RAND_50;
  reg  addresses_25_valid;
  reg [31:0] _RAND_51;
  reg [20:0] addresses_25_bits;
  reg [31:0] _RAND_52;
  reg  addresses_26_valid;
  reg [31:0] _RAND_53;
  reg [20:0] addresses_26_bits;
  reg [31:0] _RAND_54;
  reg  addresses_27_valid;
  reg [31:0] _RAND_55;
  reg [20:0] addresses_27_bits;
  reg [31:0] _RAND_56;
  reg  addresses_28_valid;
  reg [31:0] _RAND_57;
  reg [20:0] addresses_28_bits;
  reg [31:0] _RAND_58;
  reg  addresses_29_valid;
  reg [31:0] _RAND_59;
  reg [20:0] addresses_29_bits;
  reg [31:0] _RAND_60;
  reg  addresses_30_valid;
  reg [31:0] _RAND_61;
  reg [20:0] addresses_30_bits;
  reg [31:0] _RAND_62;
  reg  addresses_31_valid;
  reg [31:0] _RAND_63;
  reg [20:0] addresses_31_bits;
  reg [31:0] _RAND_64;
  reg [5:0] nextAddr;
  reg [31:0] _RAND_65;
  wire  _T_799;
  wire  _T_800;
  wire  _T_801;
  wire  _T_802;
  wire  _T_803;
  wire  _T_804;
  wire  _T_805;
  wire  _T_806;
  wire  _T_807;
  wire  _T_808;
  wire  _T_809;
  wire  _T_810;
  wire  _T_811;
  wire  _T_812;
  wire  _T_813;
  wire  _T_814;
  wire  _T_815;
  wire  _T_816;
  wire  _T_817;
  wire  _T_818;
  wire  _T_819;
  wire  _T_820;
  wire  _T_821;
  wire  _T_822;
  wire  _T_823;
  wire  _T_824;
  wire  _T_825;
  wire  _T_826;
  wire  _T_827;
  wire  _T_828;
  wire  _T_829;
  wire  _T_830;
  wire  _T_831;
  wire  _T_832;
  wire  _T_833;
  wire  _T_834;
  wire  _T_835;
  wire  _T_836;
  wire  _T_837;
  wire  _T_838;
  wire  _T_839;
  wire  _T_840;
  wire  _T_841;
  wire  _T_842;
  wire  _T_843;
  wire  _T_844;
  wire  _T_845;
  wire  _T_846;
  wire  _T_847;
  wire  _T_848;
  wire  _T_849;
  wire  _T_850;
  wire  _T_851;
  wire  _T_852;
  wire  _T_853;
  wire  _T_854;
  wire  _T_855;
  wire  _T_856;
  wire  _T_857;
  wire  _T_858;
  wire  _T_859;
  wire  _T_860;
  wire  _T_861;
  wire  _T_862;
  wire [1:0] _T_900;
  wire [1:0] _T_901;
  wire [3:0] _T_902;
  wire [1:0] _T_903;
  wire [1:0] _T_904;
  wire [3:0] _T_905;
  wire [7:0] _T_906;
  wire [1:0] _T_907;
  wire [1:0] _T_908;
  wire [3:0] _T_909;
  wire [1:0] _T_910;
  wire [1:0] _T_911;
  wire [3:0] _T_912;
  wire [7:0] _T_913;
  wire [15:0] _T_914;
  wire [1:0] _T_915;
  wire [1:0] _T_916;
  wire [3:0] _T_917;
  wire [1:0] _T_918;
  wire [1:0] _T_919;
  wire [3:0] _T_920;
  wire [7:0] _T_921;
  wire [1:0] _T_922;
  wire [1:0] _T_923;
  wire [3:0] _T_924;
  wire [1:0] _T_925;
  wire [1:0] _T_926;
  wire [3:0] _T_927;
  wire [7:0] _T_928;
  wire [15:0] _T_929;
  wire [31:0] _T_930;
  wire  _T_932;
  wire [15:0] _T_933;
  wire [15:0] _T_934;
  wire  _T_936;
  wire [15:0] _T_937;
  wire [7:0] _T_938;
  wire [7:0] _T_939;
  wire  _T_941;
  wire [7:0] _T_942;
  wire [3:0] _T_943;
  wire [3:0] _T_944;
  wire  _T_946;
  wire [3:0] _T_947;
  wire [1:0] _T_948;
  wire [1:0] _T_949;
  wire  _T_951;
  wire [1:0] _T_952;
  wire  _T_953;
  wire [1:0] _T_954;
  wire [2:0] _T_955;
  wire [3:0] _T_956;
  wire  _T_964;
  wire  _T_965;
  wire  _T_966;
  wire  _T_967;
  wire  _T_968;
  wire  _T_969;
  wire  _T_970;
  wire  _T_971;
  wire  _T_972;
  wire  _T_973;
  wire  _T_974;
  wire  _T_975;
  wire  _T_976;
  wire  _T_977;
  wire  _T_978;
  wire  _T_979;
  wire  _T_980;
  wire  _T_981;
  wire  _T_982;
  wire  _T_983;
  wire  _T_984;
  wire  _T_985;
  wire  _T_986;
  wire  _T_987;
  wire  _T_988;
  wire  _T_989;
  wire  _T_990;
  wire  _T_991;
  wire  _T_992;
  wire  _T_993;
  wire  _T_994;
  wire  _T_995;
  wire  _T_996;
  wire  _T_997;
  wire  _T_998;
  wire  _T_999;
  wire  _T_1000;
  wire  _T_1001;
  wire  _T_1002;
  wire  _T_1003;
  wire  _T_1004;
  wire  _T_1005;
  wire  _T_1006;
  wire  _T_1007;
  wire  _T_1008;
  wire  _T_1009;
  wire  _T_1010;
  wire  _T_1011;
  wire  _T_1012;
  wire  _T_1013;
  wire  _T_1014;
  wire  _T_1015;
  wire  _T_1016;
  wire  _T_1017;
  wire  _T_1018;
  wire  _T_1019;
  wire  _T_1020;
  wire  _T_1021;
  wire  _T_1022;
  wire  _T_1023;
  wire  _T_1024;
  wire  _T_1025;
  wire  _T_1026;
  wire  _T_1027;
  wire [1:0] _T_1065;
  wire [1:0] _T_1066;
  wire [3:0] _T_1067;
  wire [1:0] _T_1068;
  wire [1:0] _T_1069;
  wire [3:0] _T_1070;
  wire [7:0] _T_1071;
  wire [1:0] _T_1072;
  wire [1:0] _T_1073;
  wire [3:0] _T_1074;
  wire [1:0] _T_1075;
  wire [1:0] _T_1076;
  wire [3:0] _T_1077;
  wire [7:0] _T_1078;
  wire [15:0] _T_1079;
  wire [1:0] _T_1080;
  wire [1:0] _T_1081;
  wire [3:0] _T_1082;
  wire [1:0] _T_1083;
  wire [1:0] _T_1084;
  wire [3:0] _T_1085;
  wire [7:0] _T_1086;
  wire [1:0] _T_1087;
  wire [1:0] _T_1088;
  wire [3:0] _T_1089;
  wire [1:0] _T_1090;
  wire [1:0] _T_1091;
  wire [3:0] _T_1092;
  wire [7:0] _T_1093;
  wire [15:0] _T_1094;
  wire [31:0] _T_1095;
  wire  _T_1097;
  wire [15:0] _T_1098;
  wire [15:0] _T_1099;
  wire  _T_1101;
  wire [15:0] _T_1102;
  wire [7:0] _T_1103;
  wire [7:0] _T_1104;
  wire  _T_1106;
  wire [7:0] _T_1107;
  wire [3:0] _T_1108;
  wire [3:0] _T_1109;
  wire  _T_1111;
  wire [3:0] _T_1112;
  wire [1:0] _T_1113;
  wire [1:0] _T_1114;
  wire  _T_1116;
  wire [1:0] _T_1117;
  wire  _T_1118;
  wire [1:0] _T_1119;
  wire [2:0] _T_1120;
  wire [3:0] _T_1121;
  wire  _T_1266;
  wire [3:0] _T_1286;
  wire [6:0] _T_1297;
  wire [5:0] _T_1298;
  wire [5:0] _T_1465;
  wire  _T_1489;
  wire  _T_1490;
  wire  _T_1491;
  wire  _T_1492;
  wire  _T_1493;
  wire  _T_1494;
  wire  _T_1495;
  wire  _T_1496;
  wire  _T_1497;
  wire  _T_1498;
  wire  _T_1499;
  wire  _T_1500;
  wire  _T_1501;
  wire  _T_1502;
  wire  _T_1503;
  wire  _T_1504;
  wire  _T_1505;
  wire  _T_1506;
  wire  _T_1507;
  wire  _T_1508;
  wire  _T_1509;
  wire  _T_1510;
  wire  _T_1511;
  wire  _T_1512;
  wire  _T_1513;
  wire  _T_1514;
  wire  _T_1515;
  wire  _T_1516;
  wire  _T_1517;
  wire  _T_1518;
  wire  _T_1519;
  wire  _T_1520;
  wire  _T_1521;
  wire  _T_1522;
  wire  _T_1523;
  wire  _T_1524;
  wire  _T_1525;
  wire  _T_1526;
  wire  _T_1527;
  wire  _T_1528;
  wire  _T_1529;
  wire  _T_1530;
  wire  _T_1531;
  wire  _T_1532;
  wire  _T_1533;
  wire  _T_1534;
  wire  _T_1535;
  wire  _T_1536;
  wire  _T_1537;
  wire  _T_1538;
  wire  _T_1539;
  wire  _T_1540;
  wire  _T_1541;
  wire  _T_1542;
  wire  _T_1543;
  wire  _T_1544;
  wire  _T_1545;
  wire  _T_1546;
  wire  _T_1547;
  wire  _T_1548;
  wire  _T_1549;
  wire  _T_1550;
  wire  _T_1551;
  wire  _T_1552;
  wire [1:0] _T_1590;
  wire [1:0] _T_1591;
  wire [3:0] _T_1592;
  wire [1:0] _T_1593;
  wire [1:0] _T_1594;
  wire [3:0] _T_1595;
  wire [7:0] _T_1596;
  wire [1:0] _T_1597;
  wire [1:0] _T_1598;
  wire [3:0] _T_1599;
  wire [1:0] _T_1600;
  wire [1:0] _T_1601;
  wire [3:0] _T_1602;
  wire [7:0] _T_1603;
  wire [15:0] _T_1604;
  wire [1:0] _T_1605;
  wire [1:0] _T_1606;
  wire [3:0] _T_1607;
  wire [1:0] _T_1608;
  wire [1:0] _T_1609;
  wire [3:0] _T_1610;
  wire [7:0] _T_1611;
  wire [1:0] _T_1612;
  wire [1:0] _T_1613;
  wire [3:0] _T_1614;
  wire [1:0] _T_1615;
  wire [1:0] _T_1616;
  wire [3:0] _T_1617;
  wire [7:0] _T_1618;
  wire [15:0] _T_1619;
  wire [31:0] _T_1620;
  wire  _T_1622;
  wire [15:0] _T_1623;
  wire [15:0] _T_1624;
  wire  _T_1626;
  wire [15:0] _T_1627;
  wire [7:0] _T_1628;
  wire [7:0] _T_1629;
  wire  _T_1631;
  wire [7:0] _T_1632;
  wire [3:0] _T_1633;
  wire [3:0] _T_1634;
  wire  _T_1636;
  wire [3:0] _T_1637;
  wire [1:0] _T_1638;
  wire [1:0] _T_1639;
  wire  _T_1641;
  wire [1:0] _T_1642;
  wire  _T_1643;
  wire [1:0] _T_1644;
  wire [2:0] _T_1645;
  wire [3:0] _T_1646;
  wire [4:0] _T_1647;
  wire  _T_1649;
  wire  _T_1650;
  wire [5:0] _T_1651;
  wire  _GEN_328;
  wire  _GEN_329;
  wire  _GEN_330;
  wire  _GEN_331;
  wire  _GEN_332;
  wire  _GEN_333;
  wire  _GEN_334;
  wire  _GEN_335;
  wire  _GEN_336;
  wire  _GEN_337;
  wire  _GEN_338;
  wire  _GEN_339;
  wire  _GEN_340;
  wire  _GEN_341;
  wire  _GEN_342;
  wire  _GEN_343;
  wire  _GEN_344;
  wire  _GEN_345;
  wire  _GEN_346;
  wire  _GEN_347;
  wire  _GEN_348;
  wire  _GEN_349;
  wire  _GEN_350;
  wire  _GEN_351;
  wire  _GEN_352;
  wire  _GEN_353;
  wire  _GEN_354;
  wire  _GEN_355;
  wire  _GEN_356;
  wire  _GEN_357;
  wire  _GEN_358;
  wire  _GEN_359;
  wire [5:0] nextAddrUpdate;
  wire  _T_1675;
  wire  _T_1680;
  assign mem__T_959_addr = {_T_936,_T_956};
  assign mem__T_959_data = mem[mem__T_959_addr];
  assign mem__T_1124_addr = {_T_1101,_T_1121};
  assign mem__T_1124_data = mem[mem__T_1124_addr];
  assign mem__T_1289_addr = {_T_1266,_T_1286};
  assign mem__T_1289_data = mem[mem__T_1289_addr];
  assign mem__T_1484_data = 8'h0;
  assign mem__T_1484_addr = _T_1465[4:0];
  assign mem__T_1484_mask = 1'h0;
  assign mem__T_1484_en = 1'h0;
  assign mem__T_1670_data = io_w_1_data;
  assign mem__T_1670_addr = _T_1651[4:0];
  assign mem__T_1670_mask = io_w_1_en;
  assign mem__T_1670_en = io_w_1_en;
  assign _GEN_395 = {_T_1101,_T_1121};
  assign _GEN_404 = _T_1651[4:0];
  assign _T_799 = addresses_0_bits == io_r_0_addr;
  assign _T_800 = addresses_0_valid & _T_799;
  assign _T_801 = addresses_1_bits == io_r_0_addr;
  assign _T_802 = addresses_1_valid & _T_801;
  assign _T_803 = addresses_2_bits == io_r_0_addr;
  assign _T_804 = addresses_2_valid & _T_803;
  assign _T_805 = addresses_3_bits == io_r_0_addr;
  assign _T_806 = addresses_3_valid & _T_805;
  assign _T_807 = addresses_4_bits == io_r_0_addr;
  assign _T_808 = addresses_4_valid & _T_807;
  assign _T_809 = addresses_5_bits == io_r_0_addr;
  assign _T_810 = addresses_5_valid & _T_809;
  assign _T_811 = addresses_6_bits == io_r_0_addr;
  assign _T_812 = addresses_6_valid & _T_811;
  assign _T_813 = addresses_7_bits == io_r_0_addr;
  assign _T_814 = addresses_7_valid & _T_813;
  assign _T_815 = addresses_8_bits == io_r_0_addr;
  assign _T_816 = addresses_8_valid & _T_815;
  assign _T_817 = addresses_9_bits == io_r_0_addr;
  assign _T_818 = addresses_9_valid & _T_817;
  assign _T_819 = addresses_10_bits == io_r_0_addr;
  assign _T_820 = addresses_10_valid & _T_819;
  assign _T_821 = addresses_11_bits == io_r_0_addr;
  assign _T_822 = addresses_11_valid & _T_821;
  assign _T_823 = addresses_12_bits == io_r_0_addr;
  assign _T_824 = addresses_12_valid & _T_823;
  assign _T_825 = addresses_13_bits == io_r_0_addr;
  assign _T_826 = addresses_13_valid & _T_825;
  assign _T_827 = addresses_14_bits == io_r_0_addr;
  assign _T_828 = addresses_14_valid & _T_827;
  assign _T_829 = addresses_15_bits == io_r_0_addr;
  assign _T_830 = addresses_15_valid & _T_829;
  assign _T_831 = addresses_16_bits == io_r_0_addr;
  assign _T_832 = addresses_16_valid & _T_831;
  assign _T_833 = addresses_17_bits == io_r_0_addr;
  assign _T_834 = addresses_17_valid & _T_833;
  assign _T_835 = addresses_18_bits == io_r_0_addr;
  assign _T_836 = addresses_18_valid & _T_835;
  assign _T_837 = addresses_19_bits == io_r_0_addr;
  assign _T_838 = addresses_19_valid & _T_837;
  assign _T_839 = addresses_20_bits == io_r_0_addr;
  assign _T_840 = addresses_20_valid & _T_839;
  assign _T_841 = addresses_21_bits == io_r_0_addr;
  assign _T_842 = addresses_21_valid & _T_841;
  assign _T_843 = addresses_22_bits == io_r_0_addr;
  assign _T_844 = addresses_22_valid & _T_843;
  assign _T_845 = addresses_23_bits == io_r_0_addr;
  assign _T_846 = addresses_23_valid & _T_845;
  assign _T_847 = addresses_24_bits == io_r_0_addr;
  assign _T_848 = addresses_24_valid & _T_847;
  assign _T_849 = addresses_25_bits == io_r_0_addr;
  assign _T_850 = addresses_25_valid & _T_849;
  assign _T_851 = addresses_26_bits == io_r_0_addr;
  assign _T_852 = addresses_26_valid & _T_851;
  assign _T_853 = addresses_27_bits == io_r_0_addr;
  assign _T_854 = addresses_27_valid & _T_853;
  assign _T_855 = addresses_28_bits == io_r_0_addr;
  assign _T_856 = addresses_28_valid & _T_855;
  assign _T_857 = addresses_29_bits == io_r_0_addr;
  assign _T_858 = addresses_29_valid & _T_857;
  assign _T_859 = addresses_30_bits == io_r_0_addr;
  assign _T_860 = addresses_30_valid & _T_859;
  assign _T_861 = addresses_31_bits == io_r_0_addr;
  assign _T_862 = addresses_31_valid & _T_861;
  assign _T_900 = {_T_802,_T_800};
  assign _T_901 = {_T_806,_T_804};
  assign _T_902 = {_T_901,_T_900};
  assign _T_903 = {_T_810,_T_808};
  assign _T_904 = {_T_814,_T_812};
  assign _T_905 = {_T_904,_T_903};
  assign _T_906 = {_T_905,_T_902};
  assign _T_907 = {_T_818,_T_816};
  assign _T_908 = {_T_822,_T_820};
  assign _T_909 = {_T_908,_T_907};
  assign _T_910 = {_T_826,_T_824};
  assign _T_911 = {_T_830,_T_828};
  assign _T_912 = {_T_911,_T_910};
  assign _T_913 = {_T_912,_T_909};
  assign _T_914 = {_T_913,_T_906};
  assign _T_915 = {_T_834,_T_832};
  assign _T_916 = {_T_838,_T_836};
  assign _T_917 = {_T_916,_T_915};
  assign _T_918 = {_T_842,_T_840};
  assign _T_919 = {_T_846,_T_844};
  assign _T_920 = {_T_919,_T_918};
  assign _T_921 = {_T_920,_T_917};
  assign _T_922 = {_T_850,_T_848};
  assign _T_923 = {_T_854,_T_852};
  assign _T_924 = {_T_923,_T_922};
  assign _T_925 = {_T_858,_T_856};
  assign _T_926 = {_T_862,_T_860};
  assign _T_927 = {_T_926,_T_925};
  assign _T_928 = {_T_927,_T_924};
  assign _T_929 = {_T_928,_T_921};
  assign _T_930 = {_T_929,_T_914};
  assign _T_932 = _T_930 != 32'h0;
  assign _T_933 = _T_930[31:16];
  assign _T_934 = _T_930[15:0];
  assign _T_936 = _T_933 != 16'h0;
  assign _T_937 = _T_933 | _T_934;
  assign _T_938 = _T_937[15:8];
  assign _T_939 = _T_937[7:0];
  assign _T_941 = _T_938 != 8'h0;
  assign _T_942 = _T_938 | _T_939;
  assign _T_943 = _T_942[7:4];
  assign _T_944 = _T_942[3:0];
  assign _T_946 = _T_943 != 4'h0;
  assign _T_947 = _T_943 | _T_944;
  assign _T_948 = _T_947[3:2];
  assign _T_949 = _T_947[1:0];
  assign _T_951 = _T_948 != 2'h0;
  assign _T_952 = _T_948 | _T_949;
  assign _T_953 = _T_952[1];
  assign _T_954 = {_T_951,_T_953};
  assign _T_955 = {_T_946,_T_954};
  assign _T_956 = {_T_941,_T_955};
  assign _T_964 = addresses_0_bits == 21'h0;
  assign _T_965 = addresses_0_valid & _T_964;
  assign _T_966 = addresses_1_bits == 21'h0;
  assign _T_967 = addresses_1_valid & _T_966;
  assign _T_968 = addresses_2_bits == 21'h0;
  assign _T_969 = addresses_2_valid & _T_968;
  assign _T_970 = addresses_3_bits == 21'h0;
  assign _T_971 = addresses_3_valid & _T_970;
  assign _T_972 = addresses_4_bits == 21'h0;
  assign _T_973 = addresses_4_valid & _T_972;
  assign _T_974 = addresses_5_bits == 21'h0;
  assign _T_975 = addresses_5_valid & _T_974;
  assign _T_976 = addresses_6_bits == 21'h0;
  assign _T_977 = addresses_6_valid & _T_976;
  assign _T_978 = addresses_7_bits == 21'h0;
  assign _T_979 = addresses_7_valid & _T_978;
  assign _T_980 = addresses_8_bits == 21'h0;
  assign _T_981 = addresses_8_valid & _T_980;
  assign _T_982 = addresses_9_bits == 21'h0;
  assign _T_983 = addresses_9_valid & _T_982;
  assign _T_984 = addresses_10_bits == 21'h0;
  assign _T_985 = addresses_10_valid & _T_984;
  assign _T_986 = addresses_11_bits == 21'h0;
  assign _T_987 = addresses_11_valid & _T_986;
  assign _T_988 = addresses_12_bits == 21'h0;
  assign _T_989 = addresses_12_valid & _T_988;
  assign _T_990 = addresses_13_bits == 21'h0;
  assign _T_991 = addresses_13_valid & _T_990;
  assign _T_992 = addresses_14_bits == 21'h0;
  assign _T_993 = addresses_14_valid & _T_992;
  assign _T_994 = addresses_15_bits == 21'h0;
  assign _T_995 = addresses_15_valid & _T_994;
  assign _T_996 = addresses_16_bits == 21'h0;
  assign _T_997 = addresses_16_valid & _T_996;
  assign _T_998 = addresses_17_bits == 21'h0;
  assign _T_999 = addresses_17_valid & _T_998;
  assign _T_1000 = addresses_18_bits == 21'h0;
  assign _T_1001 = addresses_18_valid & _T_1000;
  assign _T_1002 = addresses_19_bits == 21'h0;
  assign _T_1003 = addresses_19_valid & _T_1002;
  assign _T_1004 = addresses_20_bits == 21'h0;
  assign _T_1005 = addresses_20_valid & _T_1004;
  assign _T_1006 = addresses_21_bits == 21'h0;
  assign _T_1007 = addresses_21_valid & _T_1006;
  assign _T_1008 = addresses_22_bits == 21'h0;
  assign _T_1009 = addresses_22_valid & _T_1008;
  assign _T_1010 = addresses_23_bits == 21'h0;
  assign _T_1011 = addresses_23_valid & _T_1010;
  assign _T_1012 = addresses_24_bits == 21'h0;
  assign _T_1013 = addresses_24_valid & _T_1012;
  assign _T_1014 = addresses_25_bits == 21'h0;
  assign _T_1015 = addresses_25_valid & _T_1014;
  assign _T_1016 = addresses_26_bits == 21'h0;
  assign _T_1017 = addresses_26_valid & _T_1016;
  assign _T_1018 = addresses_27_bits == 21'h0;
  assign _T_1019 = addresses_27_valid & _T_1018;
  assign _T_1020 = addresses_28_bits == 21'h0;
  assign _T_1021 = addresses_28_valid & _T_1020;
  assign _T_1022 = addresses_29_bits == 21'h0;
  assign _T_1023 = addresses_29_valid & _T_1022;
  assign _T_1024 = addresses_30_bits == 21'h0;
  assign _T_1025 = addresses_30_valid & _T_1024;
  assign _T_1026 = addresses_31_bits == 21'h0;
  assign _T_1027 = addresses_31_valid & _T_1026;
  assign _T_1065 = {_T_967,_T_965};
  assign _T_1066 = {_T_971,_T_969};
  assign _T_1067 = {_T_1066,_T_1065};
  assign _T_1068 = {_T_975,_T_973};
  assign _T_1069 = {_T_979,_T_977};
  assign _T_1070 = {_T_1069,_T_1068};
  assign _T_1071 = {_T_1070,_T_1067};
  assign _T_1072 = {_T_983,_T_981};
  assign _T_1073 = {_T_987,_T_985};
  assign _T_1074 = {_T_1073,_T_1072};
  assign _T_1075 = {_T_991,_T_989};
  assign _T_1076 = {_T_995,_T_993};
  assign _T_1077 = {_T_1076,_T_1075};
  assign _T_1078 = {_T_1077,_T_1074};
  assign _T_1079 = {_T_1078,_T_1071};
  assign _T_1080 = {_T_999,_T_997};
  assign _T_1081 = {_T_1003,_T_1001};
  assign _T_1082 = {_T_1081,_T_1080};
  assign _T_1083 = {_T_1007,_T_1005};
  assign _T_1084 = {_T_1011,_T_1009};
  assign _T_1085 = {_T_1084,_T_1083};
  assign _T_1086 = {_T_1085,_T_1082};
  assign _T_1087 = {_T_1015,_T_1013};
  assign _T_1088 = {_T_1019,_T_1017};
  assign _T_1089 = {_T_1088,_T_1087};
  assign _T_1090 = {_T_1023,_T_1021};
  assign _T_1091 = {_T_1027,_T_1025};
  assign _T_1092 = {_T_1091,_T_1090};
  assign _T_1093 = {_T_1092,_T_1089};
  assign _T_1094 = {_T_1093,_T_1086};
  assign _T_1095 = {_T_1094,_T_1079};
  assign _T_1097 = _T_1095 != 32'h0;
  assign _T_1098 = _T_1095[31:16];
  assign _T_1099 = _T_1095[15:0];
  assign _T_1101 = _T_1098 != 16'h0;
  assign _T_1102 = _T_1098 | _T_1099;
  assign _T_1103 = _T_1102[15:8];
  assign _T_1104 = _T_1102[7:0];
  assign _T_1106 = _T_1103 != 8'h0;
  assign _T_1107 = _T_1103 | _T_1104;
  assign _T_1108 = _T_1107[7:4];
  assign _T_1109 = _T_1107[3:0];
  assign _T_1111 = _T_1108 != 4'h0;
  assign _T_1112 = _T_1108 | _T_1109;
  assign _T_1113 = _T_1112[3:2];
  assign _T_1114 = _T_1112[1:0];
  assign _T_1116 = _T_1113 != 2'h0;
  assign _T_1117 = _T_1113 | _T_1114;
  assign _T_1118 = _T_1117[1];
  assign _T_1119 = {_T_1116,_T_1118};
  assign _T_1120 = {_T_1111,_T_1119};
  assign _T_1121 = {_T_1106,_T_1120};
  assign _T_1266 = _T_1098 != 16'h0;
  assign _T_1286 = {_T_1106,_T_1120};
  assign _T_1297 = nextAddr + 6'h1;
  assign _T_1298 = _T_1297[5:0];
  assign _T_1465 = _T_1097 ? {{1'd0}, _GEN_395} : nextAddr;
  assign _T_1489 = addresses_0_bits == io_w_1_addr;
  assign _T_1490 = addresses_0_valid & _T_1489;
  assign _T_1491 = addresses_1_bits == io_w_1_addr;
  assign _T_1492 = addresses_1_valid & _T_1491;
  assign _T_1493 = addresses_2_bits == io_w_1_addr;
  assign _T_1494 = addresses_2_valid & _T_1493;
  assign _T_1495 = addresses_3_bits == io_w_1_addr;
  assign _T_1496 = addresses_3_valid & _T_1495;
  assign _T_1497 = addresses_4_bits == io_w_1_addr;
  assign _T_1498 = addresses_4_valid & _T_1497;
  assign _T_1499 = addresses_5_bits == io_w_1_addr;
  assign _T_1500 = addresses_5_valid & _T_1499;
  assign _T_1501 = addresses_6_bits == io_w_1_addr;
  assign _T_1502 = addresses_6_valid & _T_1501;
  assign _T_1503 = addresses_7_bits == io_w_1_addr;
  assign _T_1504 = addresses_7_valid & _T_1503;
  assign _T_1505 = addresses_8_bits == io_w_1_addr;
  assign _T_1506 = addresses_8_valid & _T_1505;
  assign _T_1507 = addresses_9_bits == io_w_1_addr;
  assign _T_1508 = addresses_9_valid & _T_1507;
  assign _T_1509 = addresses_10_bits == io_w_1_addr;
  assign _T_1510 = addresses_10_valid & _T_1509;
  assign _T_1511 = addresses_11_bits == io_w_1_addr;
  assign _T_1512 = addresses_11_valid & _T_1511;
  assign _T_1513 = addresses_12_bits == io_w_1_addr;
  assign _T_1514 = addresses_12_valid & _T_1513;
  assign _T_1515 = addresses_13_bits == io_w_1_addr;
  assign _T_1516 = addresses_13_valid & _T_1515;
  assign _T_1517 = addresses_14_bits == io_w_1_addr;
  assign _T_1518 = addresses_14_valid & _T_1517;
  assign _T_1519 = addresses_15_bits == io_w_1_addr;
  assign _T_1520 = addresses_15_valid & _T_1519;
  assign _T_1521 = addresses_16_bits == io_w_1_addr;
  assign _T_1522 = addresses_16_valid & _T_1521;
  assign _T_1523 = addresses_17_bits == io_w_1_addr;
  assign _T_1524 = addresses_17_valid & _T_1523;
  assign _T_1525 = addresses_18_bits == io_w_1_addr;
  assign _T_1526 = addresses_18_valid & _T_1525;
  assign _T_1527 = addresses_19_bits == io_w_1_addr;
  assign _T_1528 = addresses_19_valid & _T_1527;
  assign _T_1529 = addresses_20_bits == io_w_1_addr;
  assign _T_1530 = addresses_20_valid & _T_1529;
  assign _T_1531 = addresses_21_bits == io_w_1_addr;
  assign _T_1532 = addresses_21_valid & _T_1531;
  assign _T_1533 = addresses_22_bits == io_w_1_addr;
  assign _T_1534 = addresses_22_valid & _T_1533;
  assign _T_1535 = addresses_23_bits == io_w_1_addr;
  assign _T_1536 = addresses_23_valid & _T_1535;
  assign _T_1537 = addresses_24_bits == io_w_1_addr;
  assign _T_1538 = addresses_24_valid & _T_1537;
  assign _T_1539 = addresses_25_bits == io_w_1_addr;
  assign _T_1540 = addresses_25_valid & _T_1539;
  assign _T_1541 = addresses_26_bits == io_w_1_addr;
  assign _T_1542 = addresses_26_valid & _T_1541;
  assign _T_1543 = addresses_27_bits == io_w_1_addr;
  assign _T_1544 = addresses_27_valid & _T_1543;
  assign _T_1545 = addresses_28_bits == io_w_1_addr;
  assign _T_1546 = addresses_28_valid & _T_1545;
  assign _T_1547 = addresses_29_bits == io_w_1_addr;
  assign _T_1548 = addresses_29_valid & _T_1547;
  assign _T_1549 = addresses_30_bits == io_w_1_addr;
  assign _T_1550 = addresses_30_valid & _T_1549;
  assign _T_1551 = addresses_31_bits == io_w_1_addr;
  assign _T_1552 = addresses_31_valid & _T_1551;
  assign _T_1590 = {_T_1492,_T_1490};
  assign _T_1591 = {_T_1496,_T_1494};
  assign _T_1592 = {_T_1591,_T_1590};
  assign _T_1593 = {_T_1500,_T_1498};
  assign _T_1594 = {_T_1504,_T_1502};
  assign _T_1595 = {_T_1594,_T_1593};
  assign _T_1596 = {_T_1595,_T_1592};
  assign _T_1597 = {_T_1508,_T_1506};
  assign _T_1598 = {_T_1512,_T_1510};
  assign _T_1599 = {_T_1598,_T_1597};
  assign _T_1600 = {_T_1516,_T_1514};
  assign _T_1601 = {_T_1520,_T_1518};
  assign _T_1602 = {_T_1601,_T_1600};
  assign _T_1603 = {_T_1602,_T_1599};
  assign _T_1604 = {_T_1603,_T_1596};
  assign _T_1605 = {_T_1524,_T_1522};
  assign _T_1606 = {_T_1528,_T_1526};
  assign _T_1607 = {_T_1606,_T_1605};
  assign _T_1608 = {_T_1532,_T_1530};
  assign _T_1609 = {_T_1536,_T_1534};
  assign _T_1610 = {_T_1609,_T_1608};
  assign _T_1611 = {_T_1610,_T_1607};
  assign _T_1612 = {_T_1540,_T_1538};
  assign _T_1613 = {_T_1544,_T_1542};
  assign _T_1614 = {_T_1613,_T_1612};
  assign _T_1615 = {_T_1548,_T_1546};
  assign _T_1616 = {_T_1552,_T_1550};
  assign _T_1617 = {_T_1616,_T_1615};
  assign _T_1618 = {_T_1617,_T_1614};
  assign _T_1619 = {_T_1618,_T_1611};
  assign _T_1620 = {_T_1619,_T_1604};
  assign _T_1622 = _T_1620 != 32'h0;
  assign _T_1623 = _T_1620[31:16];
  assign _T_1624 = _T_1620[15:0];
  assign _T_1626 = _T_1623 != 16'h0;
  assign _T_1627 = _T_1623 | _T_1624;
  assign _T_1628 = _T_1627[15:8];
  assign _T_1629 = _T_1627[7:0];
  assign _T_1631 = _T_1628 != 8'h0;
  assign _T_1632 = _T_1628 | _T_1629;
  assign _T_1633 = _T_1632[7:4];
  assign _T_1634 = _T_1632[3:0];
  assign _T_1636 = _T_1633 != 4'h0;
  assign _T_1637 = _T_1633 | _T_1634;
  assign _T_1638 = _T_1637[3:2];
  assign _T_1639 = _T_1637[1:0];
  assign _T_1641 = _T_1638 != 2'h0;
  assign _T_1642 = _T_1638 | _T_1639;
  assign _T_1643 = _T_1642[1];
  assign _T_1644 = {_T_1641,_T_1643};
  assign _T_1645 = {_T_1636,_T_1644};
  assign _T_1646 = {_T_1631,_T_1645};
  assign _T_1647 = {_T_1626,_T_1646};
  assign _T_1649 = _T_1622 == 1'h0;
  assign _T_1650 = io_w_1_en & _T_1649;
  assign _T_1651 = _T_1622 ? {{1'd0}, _T_1647} : nextAddr;
  assign _GEN_328 = 5'h0 == _GEN_404;
  assign _GEN_329 = 5'h1 == _GEN_404;
  assign _GEN_330 = 5'h2 == _GEN_404;
  assign _GEN_331 = 5'h3 == _GEN_404;
  assign _GEN_332 = 5'h4 == _GEN_404;
  assign _GEN_333 = 5'h5 == _GEN_404;
  assign _GEN_334 = 5'h6 == _GEN_404;
  assign _GEN_335 = 5'h7 == _GEN_404;
  assign _GEN_336 = 5'h8 == _GEN_404;
  assign _GEN_337 = 5'h9 == _GEN_404;
  assign _GEN_338 = 5'ha == _GEN_404;
  assign _GEN_339 = 5'hb == _GEN_404;
  assign _GEN_340 = 5'hc == _GEN_404;
  assign _GEN_341 = 5'hd == _GEN_404;
  assign _GEN_342 = 5'he == _GEN_404;
  assign _GEN_343 = 5'hf == _GEN_404;
  assign _GEN_344 = 5'h10 == _GEN_404;
  assign _GEN_345 = 5'h11 == _GEN_404;
  assign _GEN_346 = 5'h12 == _GEN_404;
  assign _GEN_347 = 5'h13 == _GEN_404;
  assign _GEN_348 = 5'h14 == _GEN_404;
  assign _GEN_349 = 5'h15 == _GEN_404;
  assign _GEN_350 = 5'h16 == _GEN_404;
  assign _GEN_351 = 5'h17 == _GEN_404;
  assign _GEN_352 = 5'h18 == _GEN_404;
  assign _GEN_353 = 5'h19 == _GEN_404;
  assign _GEN_354 = 5'h1a == _GEN_404;
  assign _GEN_355 = 5'h1b == _GEN_404;
  assign _GEN_356 = 5'h1c == _GEN_404;
  assign _GEN_357 = 5'h1d == _GEN_404;
  assign _GEN_358 = 5'h1e == _GEN_404;
  assign _GEN_359 = 5'h1f == _GEN_404;
  assign nextAddrUpdate = _T_1650 ? _T_1298 : nextAddr;
  assign _T_1675 = nextAddrUpdate <= 6'h20;
  assign _T_1680 = _T_1675 == 1'h0;
  assign io_r_0_data = _T_932 ? mem__T_959_data : 8'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    mem[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  addresses_0_valid = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  addresses_0_bits = _RAND_2[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  addresses_1_valid = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  addresses_1_bits = _RAND_4[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  addresses_2_valid = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  addresses_2_bits = _RAND_6[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  addresses_3_valid = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  addresses_3_bits = _RAND_8[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  addresses_4_valid = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  addresses_4_bits = _RAND_10[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  addresses_5_valid = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  addresses_5_bits = _RAND_12[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  addresses_6_valid = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  addresses_6_bits = _RAND_14[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  addresses_7_valid = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  addresses_7_bits = _RAND_16[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  addresses_8_valid = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  addresses_8_bits = _RAND_18[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  addresses_9_valid = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  addresses_9_bits = _RAND_20[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  addresses_10_valid = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  addresses_10_bits = _RAND_22[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  addresses_11_valid = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  addresses_11_bits = _RAND_24[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  addresses_12_valid = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  addresses_12_bits = _RAND_26[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  addresses_13_valid = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  addresses_13_bits = _RAND_28[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  addresses_14_valid = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  addresses_14_bits = _RAND_30[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  addresses_15_valid = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  addresses_15_bits = _RAND_32[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  addresses_16_valid = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  addresses_16_bits = _RAND_34[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  addresses_17_valid = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  addresses_17_bits = _RAND_36[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  addresses_18_valid = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  addresses_18_bits = _RAND_38[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  addresses_19_valid = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  addresses_19_bits = _RAND_40[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  addresses_20_valid = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  addresses_20_bits = _RAND_42[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  addresses_21_valid = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  addresses_21_bits = _RAND_44[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  addresses_22_valid = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  addresses_22_bits = _RAND_46[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  addresses_23_valid = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  addresses_23_bits = _RAND_48[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  addresses_24_valid = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  addresses_24_bits = _RAND_50[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  addresses_25_valid = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  addresses_25_bits = _RAND_52[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  addresses_26_valid = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  addresses_26_bits = _RAND_54[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  addresses_27_valid = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  addresses_27_bits = _RAND_56[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  addresses_28_valid = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  addresses_28_bits = _RAND_58[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  addresses_29_valid = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  addresses_29_bits = _RAND_60[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  addresses_30_valid = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  addresses_30_bits = _RAND_62[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  addresses_31_valid = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  addresses_31_bits = _RAND_64[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{$random}};
  nextAddr = _RAND_65[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(mem__T_1484_en & mem__T_1484_mask) begin
      mem[mem__T_1484_addr] <= mem__T_1484_data;
    end
    if(mem__T_1670_en & mem__T_1670_mask) begin
      mem[mem__T_1670_addr] <= mem__T_1670_data;
    end
    if (metaReset) begin
      addresses_0_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_328) begin
          addresses_0_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_0_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_328) begin
          addresses_0_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_1_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_329) begin
          addresses_1_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_1_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_329) begin
          addresses_1_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_2_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_330) begin
          addresses_2_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_2_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_330) begin
          addresses_2_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_3_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_331) begin
          addresses_3_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_3_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_331) begin
          addresses_3_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_4_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_332) begin
          addresses_4_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_4_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_332) begin
          addresses_4_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_5_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_333) begin
          addresses_5_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_5_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_333) begin
          addresses_5_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_6_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_334) begin
          addresses_6_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_6_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_334) begin
          addresses_6_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_7_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_335) begin
          addresses_7_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_7_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_335) begin
          addresses_7_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_8_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_336) begin
          addresses_8_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_8_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_336) begin
          addresses_8_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_9_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_337) begin
          addresses_9_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_9_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_337) begin
          addresses_9_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_10_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_338) begin
          addresses_10_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_10_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_338) begin
          addresses_10_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_11_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_339) begin
          addresses_11_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_11_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_339) begin
          addresses_11_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_12_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_340) begin
          addresses_12_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_12_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_340) begin
          addresses_12_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_13_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_341) begin
          addresses_13_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_13_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_341) begin
          addresses_13_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_14_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_342) begin
          addresses_14_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_14_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_342) begin
          addresses_14_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_15_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_343) begin
          addresses_15_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_15_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_343) begin
          addresses_15_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_16_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_344) begin
          addresses_16_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_16_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_344) begin
          addresses_16_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_17_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_345) begin
          addresses_17_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_17_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_345) begin
          addresses_17_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_18_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_346) begin
          addresses_18_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_18_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_346) begin
          addresses_18_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_19_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_347) begin
          addresses_19_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_19_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_347) begin
          addresses_19_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_20_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_348) begin
          addresses_20_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_20_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_348) begin
          addresses_20_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_21_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_349) begin
          addresses_21_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_21_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_349) begin
          addresses_21_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_22_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_350) begin
          addresses_22_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_22_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_350) begin
          addresses_22_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_23_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_351) begin
          addresses_23_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_23_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_351) begin
          addresses_23_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_24_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_352) begin
          addresses_24_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_24_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_352) begin
          addresses_24_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_25_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_353) begin
          addresses_25_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_25_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_353) begin
          addresses_25_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_26_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_354) begin
          addresses_26_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_26_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_354) begin
          addresses_26_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_27_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_355) begin
          addresses_27_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_27_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_355) begin
          addresses_27_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_28_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_356) begin
          addresses_28_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_28_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_356) begin
          addresses_28_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_29_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_357) begin
          addresses_29_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_29_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_357) begin
          addresses_29_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_30_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_358) begin
          addresses_30_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_30_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_358) begin
          addresses_30_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      addresses_31_valid <= 1'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_359) begin
          addresses_31_valid <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      addresses_31_bits <= 21'h0;
    end else begin
      if (io_w_1_en) begin
        if (_GEN_359) begin
          addresses_31_bits <= io_w_1_addr;
        end
      end
    end
    if (metaReset) begin
      nextAddr <= 6'h0;
    end else begin
      if (_T_1650) begin
        nextAddr <= _T_1298;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1680) begin
          $fwrite(32'h80000002,"Assertion failed: SparseMem ran out of space with size %d, increase size in ReplaceMemsTransform!\n    at SparseMem.scala:103 assert(nextAddrUpdate <= depth.U,\n",6'h20);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1680) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module SyncScratchPadMemory( // @[:Sodor3Stage.fir@3856.2]
  input         metaReset,
  input         clock, // @[:Sodor3Stage.fir@3857.4]
  input  [31:0] io_core_ports_0_req_bits_addr, // @[:Sodor3Stage.fir@3859.4]
  input  [31:0] io_core_ports_0_req_bits_data, // @[:Sodor3Stage.fir@3859.4]
  input         io_core_ports_0_req_bits_fcn, // @[:Sodor3Stage.fir@3859.4]
  input  [2:0]  io_core_ports_0_req_bits_typ, // @[:Sodor3Stage.fir@3859.4]
  output [31:0] io_core_ports_0_resp_bits_data, // @[:Sodor3Stage.fir@3859.4]
  output        _GEN_3_0,
  output        _GEN_7_0,
  output        _GEN_1_1,
  output        _GEN_4_0,
  output        _GEN_2_2,
  output        _GEN_3_4,
  output        _GEN_6_3,
  output        _GEN_0_2,
  output        _GEN_1_3,
  output        _GEN_2_4,
  output        _GEN_0_4,
  output        _GEN_5_6
);
  wire  sync_data_metaReset; // @[memory.scala 199:26:Sodor3Stage.fir@3861.4]
  wire  sync_data_clock; // @[memory.scala 199:26:Sodor3Stage.fir@3861.4]
  wire [20:0] sync_data_io_dataInstr_0_addr; // @[memory.scala 199:26:Sodor3Stage.fir@3861.4]
  wire [31:0] sync_data_io_dataInstr_0_data; // @[memory.scala 199:26:Sodor3Stage.fir@3861.4]
  wire [20:0] sync_data_io_dw_addr; // @[memory.scala 199:26:Sodor3Stage.fir@3861.4]
  wire [31:0] sync_data_io_dw_data; // @[memory.scala 199:26:Sodor3Stage.fir@3861.4]
  wire  sync_data_io_dw_en; // @[memory.scala 199:26:Sodor3Stage.fir@3861.4]
  wire  sync_data__GEN_3_0; // @[memory.scala 199:26:Sodor3Stage.fir@3861.4]
  wire  sync_data__GEN_2_2; // @[memory.scala 199:26:Sodor3Stage.fir@3861.4]
  wire  sync_data__GEN_1_3; // @[memory.scala 199:26:Sodor3Stage.fir@3861.4]
  wire  sync_data__GEN_0_4; // @[memory.scala 199:26:Sodor3Stage.fir@3861.4]
  reg [2:0] req_typi; // @[memory.scala 213:22:Sodor3Stage.fir@3883.4]
  reg [31:0] _RAND_0;
  wire  _T_233; // @[memory.scala 218:17:Sodor3Stage.fir@3885.4]
  wire  _T_234; // @[memory.scala 218:52:Sodor3Stage.fir@3886.4]
  wire [23:0] _T_238; // @[Bitwise.scala 72:12:Sodor3Stage.fir@3888.4]
  wire [7:0] _T_239; // @[memory.scala 218:67:Sodor3Stage.fir@3889.4]
  wire [31:0] _T_240; // @[Cat.scala 30:58:Sodor3Stage.fir@3890.4]
  wire  _T_241; // @[memory.scala 219:17:Sodor3Stage.fir@3891.4]
  wire  _T_242; // @[memory.scala 219:52:Sodor3Stage.fir@3892.4]
  wire [15:0] _T_246; // @[Bitwise.scala 72:12:Sodor3Stage.fir@3894.4]
  wire [15:0] _T_247; // @[memory.scala 219:68:Sodor3Stage.fir@3895.4]
  wire [31:0] _T_248; // @[Cat.scala 30:58:Sodor3Stage.fir@3896.4]
  wire  _T_249; // @[memory.scala 220:17:Sodor3Stage.fir@3897.4]
  wire [31:0] _T_256; // @[Cat.scala 30:58:Sodor3Stage.fir@3900.4]
  wire  _T_257; // @[memory.scala 221:17:Sodor3Stage.fir@3901.4]
  wire [31:0] _T_264; // @[Cat.scala 30:58:Sodor3Stage.fir@3904.4]
  wire [31:0] _T_265; // @[Mux.scala 61:16:Sodor3Stage.fir@3905.4]
  wire [31:0] _T_266; // @[Mux.scala 61:16:Sodor3Stage.fir@3906.4]
  wire [31:0] _T_267; // @[Mux.scala 61:16:Sodor3Stage.fir@3907.4]
  wire [1:0] _T_275; // @[memory.scala 227:79:Sodor3Stage.fir@3916.6]
  wire [4:0] _GEN_8; // @[memory.scala 227:85:Sodor3Stage.fir@3917.6]
  wire [4:0] _T_276; // @[memory.scala 227:85:Sodor3Stage.fir@3917.6]
  wire [62:0] _GEN_10; // @[memory.scala 227:66:Sodor3Stage.fir@3918.6]
  wire [62:0] _T_277; // @[memory.scala 227:66:Sodor3Stage.fir@3918.6]
  wire [29:0] _T_278; // @[memory.scala 228:44:Sodor3Stage.fir@3920.6]
  wire [31:0] _T_280; // @[Cat.scala 30:58:Sodor3Stage.fir@3921.6]
  SyncMem sync_data ( // @[memory.scala 199:26:Sodor3Stage.fir@3861.4]
    .metaReset(sync_data_metaReset),
    .clock(sync_data_clock),
    .io_dataInstr_0_addr(sync_data_io_dataInstr_0_addr),
    .io_dataInstr_0_data(sync_data_io_dataInstr_0_data),
    .io_dw_addr(sync_data_io_dw_addr),
    .io_dw_data(sync_data_io_dw_data),
    .io_dw_en(sync_data_io_dw_en),
    ._GEN_3_0(sync_data__GEN_3_0),
    ._GEN_2_2(sync_data__GEN_2_2),
    ._GEN_1_3(sync_data__GEN_1_3),
    ._GEN_0_4(sync_data__GEN_0_4)
  );
  assign sync_data_metaReset = metaReset;
  assign _T_233 = req_typi == 3'h1; // @[memory.scala 218:17:Sodor3Stage.fir@3885.4]
  assign _T_234 = sync_data_io_dataInstr_0_data[7]; // @[memory.scala 218:52:Sodor3Stage.fir@3886.4]
  assign _T_238 = _T_234 ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12:Sodor3Stage.fir@3888.4]
  assign _T_239 = sync_data_io_dataInstr_0_data[7:0]; // @[memory.scala 218:67:Sodor3Stage.fir@3889.4]
  assign _T_240 = {_T_238,_T_239}; // @[Cat.scala 30:58:Sodor3Stage.fir@3890.4]
  assign _T_241 = req_typi == 3'h2; // @[memory.scala 219:17:Sodor3Stage.fir@3891.4]
  assign _T_242 = sync_data_io_dataInstr_0_data[15]; // @[memory.scala 219:52:Sodor3Stage.fir@3892.4]
  assign _T_246 = _T_242 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:Sodor3Stage.fir@3894.4]
  assign _T_247 = sync_data_io_dataInstr_0_data[15:0]; // @[memory.scala 219:68:Sodor3Stage.fir@3895.4]
  assign _T_248 = {_T_246,_T_247}; // @[Cat.scala 30:58:Sodor3Stage.fir@3896.4]
  assign _T_249 = req_typi == 3'h5; // @[memory.scala 220:17:Sodor3Stage.fir@3897.4]
  assign _T_256 = {24'h0,_T_239}; // @[Cat.scala 30:58:Sodor3Stage.fir@3900.4]
  assign _T_257 = req_typi == 3'h6; // @[memory.scala 221:17:Sodor3Stage.fir@3901.4]
  assign _T_264 = {16'h0,_T_247}; // @[Cat.scala 30:58:Sodor3Stage.fir@3904.4]
  assign _T_265 = _T_257 ? _T_264 : sync_data_io_dataInstr_0_data; // @[Mux.scala 61:16:Sodor3Stage.fir@3905.4]
  assign _T_266 = _T_249 ? _T_256 : _T_265; // @[Mux.scala 61:16:Sodor3Stage.fir@3906.4]
  assign _T_267 = _T_241 ? _T_248 : _T_266; // @[Mux.scala 61:16:Sodor3Stage.fir@3907.4]
  assign _T_275 = io_core_ports_0_req_bits_addr[1:0]; // @[memory.scala 227:79:Sodor3Stage.fir@3916.6]
  assign _GEN_8 = {{3'd0}, _T_275}; // @[memory.scala 227:85:Sodor3Stage.fir@3917.6]
  assign _T_276 = _GEN_8 << 3; // @[memory.scala 227:85:Sodor3Stage.fir@3917.6]
  assign _GEN_10 = {{31'd0}, io_core_ports_0_req_bits_data}; // @[memory.scala 227:66:Sodor3Stage.fir@3918.6]
  assign _T_277 = _GEN_10 << _T_276; // @[memory.scala 227:66:Sodor3Stage.fir@3918.6]
  assign _T_278 = io_core_ports_0_req_bits_addr[31:2]; // @[memory.scala 228:44:Sodor3Stage.fir@3920.6]
  assign _T_280 = {_T_278,2'h0}; // @[Cat.scala 30:58:Sodor3Stage.fir@3921.6]
  assign io_core_ports_0_resp_bits_data = _T_233 ? _T_240 : _T_267;
  assign _GEN_3_0 = sync_data__GEN_3_0;
  assign _GEN_7_0 = req_typi == 3'h1;
  assign _GEN_1_1 = sync_data_io_dataInstr_0_data[15];
  assign _GEN_4_0 = req_typi == 3'h2;
  assign _GEN_2_2 = sync_data__GEN_2_2;
  assign _GEN_3_4 = req_typi == 3'h5;
  assign _GEN_6_3 = io_core_ports_0_req_bits_typ == 3'h1;
  assign _GEN_0_2 = sync_data_io_dataInstr_0_data[7];
  assign _GEN_1_3 = sync_data__GEN_1_3;
  assign _GEN_2_4 = req_typi == 3'h6;
  assign _GEN_0_4 = sync_data__GEN_0_4;
  assign _GEN_5_6 = io_core_ports_0_req_bits_typ == 3'h2;
  assign sync_data_clock = clock;
  assign sync_data_io_dataInstr_0_addr = io_core_ports_0_req_bits_addr[20:0];
  assign sync_data_io_dw_addr = _T_280[20:0];
  assign sync_data_io_dw_data = _T_277[31:0];
  assign sync_data_io_dw_en = io_core_ports_0_req_bits_fcn;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  req_typi = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (metaReset) begin
      req_typi <= 3'h0;
    end else begin
      req_typi <= io_core_ports_0_req_bits_typ;
    end
  end
endmodule
